module database(clk,datata,re,address,we,dp,address_p);

parameter SIZE=0;

input clk;
output reg signed [SIZE-1:0] datata;
input re,we;
input [12:0] address;
input signed [SIZE-1:0] dp;
input [12:0] address_p;

reg signed [SIZE-1:0] storage [5459:0];

initial begin

storage[0] =  11'b0;
storage[1] =  11'b0;
storage[2] =  11'b0;
storage[3] =  11'b0;
storage[4] =  11'b0;
storage[5] =  11'b0;
storage[6] =  11'b0;
storage[7] =  11'b0;
storage[8] =  11'b0;
storage[9] =  11'b0;
storage[10] =  11'b0;
storage[11] =  11'b0;
storage[12] =  11'b0;
storage[13] =  11'b0;
storage[14] =  11'b0;
storage[15] =  11'b0;
storage[16] =  11'b0;
storage[17] =  11'b0;
storage[18] =  11'b0;
storage[19] =  11'b0;
storage[20] =  11'b0;
storage[21] =  11'b0;
storage[22] =  11'b0;
storage[23] =  11'b0;
storage[24] =  11'b0;
storage[25] =  11'b0;
storage[26] =  11'b0;
storage[27] =  11'b0;
storage[28] =  11'b0;
storage[29] =  11'b0;
storage[30] =  11'b0;
storage[31] =  11'b0;
storage[32] =  11'b0;
storage[33] =  11'b0;
storage[34] =  11'b0;
storage[35] =  11'b0;
storage[36] =  11'b0;
storage[37] =  11'b0;
storage[38] =  11'b0;
storage[39] =  11'b0;
storage[40] =  11'b0;
storage[41] =  11'b0;
storage[42] =  11'b0;
storage[43] =  11'b0;
storage[44] =  11'b0;
storage[45] =  11'b0;
storage[46] =  11'b0;
storage[47] =  11'b0;
storage[48] =  11'b0;
storage[49] =  11'b0;
storage[50] =  11'b0;
storage[51] =  11'b0;
storage[52] =  11'b0;
storage[53] =  11'b0;
storage[54] =  11'b0;
storage[55] =  11'b0;
storage[56] =  11'b0;
storage[57] =  11'b0;
storage[58] =  11'b0;
storage[59] =  11'b0;
storage[60] =  11'b0;
storage[61] =  11'b0;
storage[62] =  11'b0;
storage[63] =  11'b0;
storage[64] =  11'b0;
storage[65] =  11'b0;
storage[66] =  11'b0;
storage[67] =  11'b0;
storage[68] =  11'b0;
storage[69] =  11'b0;
storage[70] =  11'b0;
storage[71] =  11'b0;
storage[72] =  11'b0;
storage[73] =  11'b0;
storage[74] =  11'b0;
storage[75] =  11'b0;
storage[76] =  11'b0;
storage[77] =  11'b0;
storage[78] =  11'b0;
storage[79] =  11'b0;
storage[80] =  11'b0;
storage[81] =  11'b0;
storage[82] =  11'b0;
storage[83] =  11'b0;
storage[84] =  11'b0;
storage[85] =  11'b0;
storage[86] =  11'b0;
storage[87] =  11'b0;
storage[88] =  11'b0;
storage[89] =  11'b0;
storage[90] =  11'b0;
storage[91] =  11'b0;
storage[92] =  11'b0;
storage[93] =  11'b0;
storage[94] =  11'b0;
storage[95] =  11'b0;
storage[96] =  11'b0;
storage[97] =  11'b0;
storage[98] =  11'b0;
storage[99] =  11'b0;
storage[100] =  11'b0;
storage[101] =  11'b0;
storage[102] =  11'b0;
storage[103] =  11'b0;
storage[104] =  11'b0;
storage[105] =  11'b0;
storage[106] =  11'b0;
storage[107] =  11'b0;
storage[108] =  11'b0;
storage[109] =  11'b0;
storage[110] =  11'b0;
storage[111] =  11'b0;
storage[112] =  11'b0;
storage[113] =  11'b0;
storage[114] =  11'b0;
storage[115] =  11'b0;
storage[116] =  11'b0;
storage[117] =  11'b0;
storage[118] =  11'b0;
storage[119] =  11'b0;
storage[120] =  11'b0;
storage[121] =  11'b0;
storage[122] =  11'b0;
storage[123] =  11'b0;
storage[124] =  11'b0;
storage[125] =  11'b0;
storage[126] =  11'b0;
storage[127] =  11'b0;
storage[128] =  11'b0;
storage[129] =  11'b0;
storage[130] =  11'b0;
storage[131] =  11'b0;
storage[132] =  11'b0;
storage[133] =  11'b0;
storage[134] =  11'b0;
storage[135] =  11'b0;
storage[136] =  11'b0;
storage[137] =  11'b0;
storage[138] =  11'b0;
storage[139] =  11'b0;
storage[140] =  11'b0;
storage[141] =  11'b0;
storage[142] =  11'b0;
storage[143] =  11'b0;
storage[144] =  11'b0;
storage[145] =  11'b0;
storage[146] =  11'b0;
storage[147] =  11'b0;
storage[148] =  11'b0;
storage[149] =  11'b0;
storage[150] =  11'b0;
storage[151] =  11'b0;
storage[152] =  11'b0;
storage[153] =  11'b0;
storage[154] =  11'b0;
storage[155] =  11'b0;
storage[156] =  11'b0;
storage[157] =  11'b0;
storage[158] =  11'b0;
storage[159] =  11'b0;
storage[160] =  11'b0;
storage[161] =  11'b0;
storage[162] =  11'b0;
storage[163] =  11'b0;
storage[164] =  11'b0;
storage[165] =  11'b0;
storage[166] =  11'b0;
storage[167] =  11'b0;
storage[168] =  11'b0;
storage[169] =  11'b0;
storage[170] =  11'b0;
storage[171] =  11'b0;
storage[172] =  11'b0;
storage[173] =  11'b0;
storage[174] =  11'b0;
storage[175] =  11'b0;
storage[176] =  11'b0;
storage[177] =  11'b0;
storage[178] =  11'b0;
storage[179] =  11'b0;
storage[180] =  11'b0;
storage[181] =  11'b0;
storage[182] =  11'b0;
storage[183] =  11'b0;
storage[184] =  11'b0;
storage[185] =  11'b0;
storage[186] =  11'b0;
storage[187] =  11'b0;
storage[188] =  11'b0;
storage[189] =  11'b0;
storage[190] =  11'b0;
storage[191] =  11'b0;
storage[192] =  11'b0;
storage[193] =  11'b0;
storage[194] =  11'b0;
storage[195] =  11'b0;
storage[196] =  11'b0;
storage[197] =  11'b0;
storage[198] =  11'b0;
storage[199] =  11'b0;
storage[200] =  11'b0;
storage[201] =  11'b0;
storage[202] =  11'b0;
storage[203] =  11'b0;
storage[204] =  11'b0;
storage[205] =  11'b0;
storage[206] =  11'b0;
storage[207] =  11'b0;
storage[208] =  11'b0;
storage[209] =  11'b0;
storage[210] =  11'b0;
storage[211] =  11'b0;
storage[212] =  11'b0;
storage[213] =  11'b0;
storage[214] =  11'b0;
storage[215] =  11'b0;
storage[216] =  11'b0;
storage[217] =  11'b0;
storage[218] =  11'b0;
storage[219] =  11'b0;
storage[220] =  11'b0;
storage[221] =  11'b0;
storage[222] =  11'b0;
storage[223] =  11'b0;
storage[224] =  11'b0;
storage[225] =  11'b0;
storage[226] =  11'b0;
storage[227] =  11'b0;
storage[228] =  11'b0;
storage[229] =  11'b0;
storage[230] =  11'b0;
storage[231] =  11'b0;
storage[232] =  11'b0;
storage[233] =  11'b0;
storage[234] =  11'b0;
storage[235] =  11'b0;
storage[236] =  11'b0;
storage[237] =  11'b0;
storage[238] =  11'b0;
storage[239] =  11'b0;
storage[240] =  11'b0;
storage[241] =  11'b0;
storage[242] =  11'b0;
storage[243] =  11'b0;
storage[244] =  11'b0;
storage[245] =  11'b0;
storage[246] =  11'b0;
storage[247] =  11'b0;
storage[248] =  11'b0;
storage[249] =  11'b0;
storage[250] =  11'b0;
storage[251] =  11'b0;
storage[252] =  11'b0;
storage[253] =  11'b0;
storage[254] =  11'b0;
storage[255] =  11'b0;
storage[256] =  11'b0;
storage[257] =  11'b0;
storage[258] =  11'b0;
storage[259] =  11'b0;
storage[260] =  11'b0;
storage[261] =  11'b0;
storage[262] =  11'b0;
storage[263] =  11'b0;
storage[264] =  11'b0;
storage[265] =  11'b0;
storage[266] =  11'b0;
storage[267] =  11'b0;
storage[268] =  11'b0;
storage[269] =  11'b0;
storage[270] =  11'b0;
storage[271] =  11'b0;
storage[272] =  11'b0;
storage[273] =  11'b0;
storage[274] =  11'b0;
storage[275] =  11'b0;
storage[276] =  11'b0;
storage[277] =  11'b0;
storage[278] =  11'b0;
storage[279] =  11'b0;
storage[280] =  11'b0;
storage[281] =  11'b0;
storage[282] =  11'b0;
storage[283] =  11'b0;
storage[284] =  11'b0;
storage[285] =  11'b0;
storage[286] =  11'b0;
storage[287] =  11'b0;
storage[288] =  11'b0;
storage[289] =  11'b0;
storage[290] =  11'b0;
storage[291] =  11'b0;
storage[292] =  11'b0;
storage[293] =  11'b0;
storage[294] =  11'b0;
storage[295] =  11'b0;
storage[296] =  11'b0;
storage[297] =  11'b0;
storage[298] =  11'b0;
storage[299] =  11'b0;
storage[300] =  11'b0;
storage[301] =  11'b0;
storage[302] =  11'b0;
storage[303] =  11'b0;
storage[304] =  11'b0;
storage[305] =  11'b0;
storage[306] =  11'b0;
storage[307] =  11'b0;
storage[308] =  11'b0;
storage[309] =  11'b0;
storage[310] =  11'b0;
storage[311] =  11'b0;
storage[312] =  11'b0;
storage[313] =  11'b0;
storage[314] =  11'b0;
storage[315] =  11'b0;
storage[316] =  11'b0;
storage[317] =  11'b0;
storage[318] =  11'b0;
storage[319] =  11'b0;
storage[320] =  11'b0;
storage[321] =  11'b0;
storage[322] =  11'b0;
storage[323] =  11'b0;
storage[324] =  11'b0;
storage[325] =  11'b0;
storage[326] =  11'b0;
storage[327] =  11'b0;
storage[328] =  11'b0;
storage[329] =  11'b0;
storage[330] =  11'b0;
storage[331] =  11'b0;
storage[332] =  11'b0;
storage[333] =  11'b0;
storage[334] =  11'b0;
storage[335] =  11'b0;
storage[336] =  11'b0;
storage[337] =  11'b0;
storage[338] =  11'b0;
storage[339] =  11'b0;
storage[340] =  11'b0;
storage[341] =  11'b0;
storage[342] =  11'b0;
storage[343] =  11'b0;
storage[344] =  11'b0;
storage[345] =  11'b0;
storage[346] =  11'b0;
storage[347] =  11'b0;
storage[348] =  11'b0;
storage[349] =  11'b0;
storage[350] =  11'b0;
storage[351] =  11'b0;
storage[352] =  11'b0;
storage[353] =  11'b0;
storage[354] =  11'b0;
storage[355] =  11'b0;
storage[356] =  11'b0;
storage[357] =  11'b0;
storage[358] =  11'b0;
storage[359] =  11'b0;
storage[360] =  11'b0;
storage[361] =  11'b0;
storage[362] =  11'b0;
storage[363] =  11'b0;
storage[364] =  11'b0;
storage[365] =  11'b0;
storage[366] =  11'b0;
storage[367] =  11'b0;
storage[368] =  11'b0;
storage[369] =  11'b0;
storage[370] =  11'b0;
storage[371] =  11'b0;
storage[372] =  11'b0;
storage[373] =  11'b0;
storage[374] =  11'b0;
storage[375] =  11'b0;
storage[376] =  11'b0;
storage[377] =  11'b0;
storage[378] =  11'b0;
storage[379] =  11'b0;
storage[380] =  11'b0;
storage[381] =  11'b0;
storage[382] =  11'b0;
storage[383] =  11'b0;
storage[384] =  11'b0;
storage[385] =  11'b0;
storage[386] =  11'b0;
storage[387] =  11'b0;
storage[388] =  11'b0;
storage[389] =  11'b0;
storage[390] =  11'b0;
storage[391] =  11'b0;
storage[392] =  11'b0;
storage[393] =  11'b0;
storage[394] =  11'b0;
storage[395] =  11'b0;
storage[396] =  11'b0;
storage[397] =  11'b0;
storage[398] =  11'b0;
storage[399] =  11'b0;
storage[400] =  11'b0;
storage[401] =  11'b0;
storage[402] =  11'b0;
storage[403] =  11'b0;
storage[404] =  11'b0;
storage[405] =  11'b0;
storage[406] =  11'b0;
storage[407] =  11'b0;
storage[408] =  11'b0;
storage[409] =  11'b0;
storage[410] =  11'b0;
storage[411] =  11'b0;
storage[412] =  11'b0;
storage[413] =  11'b0;
storage[414] =  11'b0;
storage[415] =  11'b0;
storage[416] =  11'b0;
storage[417] =  11'b0;
storage[418] =  11'b0;
storage[419] =  11'b0;
storage[420] =  11'b0;
storage[421] =  11'b0;
storage[422] =  11'b0;
storage[423] =  11'b0;
storage[424] =  11'b0;
storage[425] =  11'b0;
storage[426] =  11'b0;
storage[427] =  11'b0;
storage[428] =  11'b0;
storage[429] =  11'b0;
storage[430] =  11'b0;
storage[431] =  11'b0;
storage[432] =  11'b0;
storage[433] =  11'b0;
storage[434] =  11'b0;
storage[435] =  11'b0;
storage[436] =  11'b0;
storage[437] =  11'b0;
storage[438] =  11'b0;
storage[439] =  11'b0;
storage[440] =  11'b0;
storage[441] =  11'b0;
storage[442] =  11'b0;
storage[443] =  11'b0;
storage[444] =  11'b0;
storage[445] =  11'b0;
storage[446] =  11'b0;
storage[447] =  11'b0;
storage[448] =  11'b0;
storage[449] =  11'b0;
storage[450] =  11'b0;
storage[451] =  11'b0;
storage[452] =  11'b0;
storage[453] =  11'b0;
storage[454] =  11'b0;
storage[455] =  11'b0;
storage[456] =  11'b0;
storage[457] =  11'b0;
storage[458] =  11'b0;
storage[459] =  11'b0;
storage[460] =  11'b0;
storage[461] =  11'b0;
storage[462] =  11'b0;
storage[463] =  11'b0;
storage[464] =  11'b0;
storage[465] =  11'b0;
storage[466] =  11'b0;
storage[467] =  11'b0;
storage[468] =  11'b0;
storage[469] =  11'b0;
storage[470] =  11'b0;
storage[471] =  11'b0;
storage[472] =  11'b0;
storage[473] =  11'b0;
storage[474] =  11'b0;
storage[475] =  11'b0;
storage[476] =  11'b0;
storage[477] =  11'b0;
storage[478] =  11'b0;
storage[479] =  11'b0;
storage[480] =  11'b0;
storage[481] =  11'b0;
storage[482] =  11'b0;
storage[483] =  11'b0;
storage[484] =  11'b0;
storage[485] =  11'b0;
storage[486] =  11'b0;
storage[487] =  11'b0;
storage[488] =  11'b0;
storage[489] =  11'b0;
storage[490] =  11'b0;
storage[491] =  11'b0;
storage[492] =  11'b0;
storage[493] =  11'b0;
storage[494] =  11'b0;
storage[495] =  11'b0;
storage[496] =  11'b0;
storage[497] =  11'b0;
storage[498] =  11'b0;
storage[499] =  11'b0;
storage[500] =  11'b0;
storage[501] =  11'b0;
storage[502] =  11'b0;
storage[503] =  11'b0;
storage[504] =  11'b0;
storage[505] =  11'b0;
storage[506] =  11'b0;
storage[507] =  11'b0;
storage[508] =  11'b0;
storage[509] =  11'b0;
storage[510] =  11'b0;
storage[511] =  11'b0;
storage[512] =  11'b0;
storage[513] =  11'b0;
storage[514] =  11'b0;
storage[515] =  11'b0;
storage[516] =  11'b0;
storage[517] =  11'b0;
storage[518] =  11'b0;
storage[519] =  11'b0;
storage[520] =  11'b0;
storage[521] =  11'b0;
storage[522] =  11'b0;
storage[523] =  11'b0;
storage[524] =  11'b0;
storage[525] =  11'b0;
storage[526] =  11'b0;
storage[527] =  11'b0;
storage[528] =  11'b0;
storage[529] =  11'b0;
storage[530] =  11'b0;
storage[531] =  11'b0;
storage[532] =  11'b0;
storage[533] =  11'b0;
storage[534] =  11'b0;
storage[535] =  11'b0;
storage[536] =  11'b0;
storage[537] =  11'b0;
storage[538] =  11'b0;
storage[539] =  11'b0;
storage[540] =  11'b0;
storage[541] =  11'b0;
storage[542] =  11'b0;
storage[543] =  11'b0;
storage[544] =  11'b0;
storage[545] =  11'b0;
storage[546] =  11'b0;
storage[547] =  11'b0;
storage[548] =  11'b0;
storage[549] =  11'b0;
storage[550] =  11'b0;
storage[551] =  11'b0;
storage[552] =  11'b0;
storage[553] =  11'b0;
storage[554] =  11'b0;
storage[555] =  11'b0;
storage[556] =  11'b0;
storage[557] =  11'b0;
storage[558] =  11'b0;
storage[559] =  11'b0;
storage[560] =  11'b0;
storage[561] =  11'b0;
storage[562] =  11'b0;
storage[563] =  11'b0;
storage[564] =  11'b0;
storage[565] =  11'b0;
storage[566] =  11'b0;
storage[567] =  11'b0;
storage[568] =  11'b0;
storage[569] =  11'b0;
storage[570] =  11'b0;
storage[571] =  11'b0;
storage[572] =  11'b0;
storage[573] =  11'b0;
storage[574] =  11'b0;
storage[575] =  11'b0;
storage[576] =  11'b0;
storage[577] =  11'b0;
storage[578] =  11'b0;
storage[579] =  11'b0;
storage[580] =  11'b0;
storage[581] =  11'b0;
storage[582] =  11'b0;
storage[583] =  11'b0;
storage[584] =  11'b0;
storage[585] =  11'b0;
storage[586] =  11'b0;
storage[587] =  11'b0;
storage[588] =  11'b0;
storage[589] =  11'b0;
storage[590] =  11'b0;
storage[591] =  11'b0;
storage[592] =  11'b0;
storage[593] =  11'b0;
storage[594] =  11'b0;
storage[595] =  11'b0;
storage[596] =  11'b0;
storage[597] =  11'b0;
storage[598] =  11'b0;
storage[599] =  11'b0;
storage[600] =  11'b0;
storage[601] =  11'b0;
storage[602] =  11'b0;
storage[603] =  11'b0;
storage[604] =  11'b0;
storage[605] =  11'b0;
storage[606] =  11'b0;
storage[607] =  11'b0;
storage[608] =  11'b0;
storage[609] =  11'b0;
storage[610] =  11'b0;
storage[611] =  11'b0;
storage[612] =  11'b0;
storage[613] =  11'b0;
storage[614] =  11'b0;
storage[615] =  11'b0;
storage[616] =  11'b0;
storage[617] =  11'b0;
storage[618] =  11'b0;
storage[619] =  11'b0;
storage[620] =  11'b0;
storage[621] =  11'b0;
storage[622] =  11'b0;
storage[623] =  11'b0;
storage[624] =  11'b0;
storage[625] =  11'b0;
storage[626] =  11'b0;
storage[627] =  11'b0;
storage[628] =  11'b0;
storage[629] =  11'b0;
storage[630] =  11'b0;
storage[631] =  11'b0;
storage[632] =  11'b0;
storage[633] =  11'b0;
storage[634] =  11'b0;
storage[635] =  11'b0;
storage[636] =  11'b0;
storage[637] =  11'b0;
storage[638] =  11'b0;
storage[639] =  11'b0;
storage[640] =  11'b0;
storage[641] =  11'b0;
storage[642] =  11'b0;
storage[643] =  11'b0;
storage[644] =  11'b0;
storage[645] =  11'b0;
storage[646] =  11'b0;
storage[647] =  11'b0;
storage[648] =  11'b0;
storage[649] =  11'b0;
storage[650] =  11'b0;
storage[651] =  11'b0;
storage[652] =  11'b0;
storage[653] =  11'b0;
storage[654] =  11'b0;
storage[655] =  11'b0;
storage[656] =  11'b0;
storage[657] =  11'b0;
storage[658] =  11'b0;
storage[659] =  11'b0;
storage[660] =  11'b0;
storage[661] =  11'b0;
storage[662] =  11'b0;
storage[663] =  11'b0;
storage[664] =  11'b0;
storage[665] =  11'b0;
storage[666] =  11'b0;
storage[667] =  11'b0;
storage[668] =  11'b0;
storage[669] =  11'b0;
storage[670] =  11'b0;
storage[671] =  11'b0;
storage[672] =  11'b0;
storage[673] =  11'b0;
storage[674] =  11'b0;
storage[675] =  11'b0;
storage[676] =  11'b0;
storage[677] =  11'b0;
storage[678] =  11'b0;
storage[679] =  11'b0;
storage[680] =  11'b0;
storage[681] =  11'b0;
storage[682] =  11'b0;
storage[683] =  11'b0;
storage[684] =  11'b0;
storage[685] =  11'b0;
storage[686] =  11'b0;
storage[687] =  11'b0;
storage[688] =  11'b0;
storage[689] =  11'b0;
storage[690] =  11'b0;
storage[691] =  11'b0;
storage[692] =  11'b0;
storage[693] =  11'b0;
storage[694] =  11'b0;
storage[695] =  11'b0;
storage[696] =  11'b0;
storage[697] =  11'b0;
storage[698] =  11'b0;
storage[699] =  11'b0;
storage[700] =  11'b0;
storage[701] =  11'b0;
storage[702] =  11'b0;
storage[703] =  11'b0;
storage[704] =  11'b0;
storage[705] =  11'b0;
storage[706] =  11'b0;
storage[707] =  11'b0;
storage[708] =  11'b0;
storage[709] =  11'b0;
storage[710] =  11'b0;
storage[711] =  11'b0;
storage[712] =  11'b0;
storage[713] =  11'b0;
storage[714] =  11'b0;
storage[715] =  11'b0;
storage[716] =  11'b0;
storage[717] =  11'b0;
storage[718] =  11'b0;
storage[719] =  11'b0;
storage[720] =  11'b0;
storage[721] =  11'b0;
storage[722] =  11'b0;
storage[723] =  11'b0;
storage[724] =  11'b0;
storage[725] =  11'b0;
storage[726] =  11'b0;
storage[727] =  11'b0;
storage[728] =  11'b0;
storage[729] =  11'b0;
storage[730] =  11'b0;
storage[731] =  11'b0;
storage[732] =  11'b0;
storage[733] =  11'b0;
storage[734] =  11'b0;
storage[735] =  11'b0;
storage[736] =  11'b0;
storage[737] =  11'b0;
storage[738] =  11'b0;
storage[739] =  11'b0;
storage[740] =  11'b0;
storage[741] =  11'b0;
storage[742] =  11'b0;
storage[743] =  11'b0;
storage[744] =  11'b0;
storage[745] =  11'b0;
storage[746] =  11'b0;
storage[747] =  11'b0;
storage[748] =  11'b0;
storage[749] =  11'b0;
storage[750] =  11'b0;
storage[751] =  11'b0;
storage[752] =  11'b0;
storage[753] =  11'b0;
storage[754] =  11'b0;
storage[755] =  11'b0;
storage[756] =  11'b0;
storage[757] =  11'b0;
storage[758] =  11'b0;
storage[759] =  11'b0;
storage[760] =  11'b0;
storage[761] =  11'b0;
storage[762] =  11'b0;
storage[763] =  11'b0;
storage[764] =  11'b0;
storage[765] =  11'b0;
storage[766] =  11'b0;
storage[767] =  11'b0;
storage[768] =  11'b0;
storage[769] =  11'b0;
storage[770] =  11'b0;
storage[771] =  11'b0;
storage[772] =  11'b0;
storage[773] =  11'b0;
storage[774] =  11'b0;
storage[775] =  11'b0;
storage[776] =  11'b0;
storage[777] =  11'b0;
storage[778] =  11'b0;
storage[779] =  11'b0;
storage[780] =  11'b0;
storage[781] =  11'b0;
storage[782] =  11'b0;
storage[783] =  11'b0;
storage[784] =  11'b00000011111; // 31
storage[785] =  11'b00010101101; // 173
storage[786] = -11'b00001101100; // -108
storage[787] =  11'b00100011100; // 284
storage[788] = -11'b00001111110; // -126
storage[789] = -11'b00001000111; // -71
storage[790] = -11'b00000111110; // -62
storage[791] = -11'b00000001101; // -13
storage[792] = -11'b00000110011; // -51
storage[793] = -11'b00010001110; // -142
storage[794] = -11'b00010001010; // -138
storage[795] = -11'b00010111100; // -188
storage[796] =  11'b00001111111; // 127
storage[797] =  11'b00011000000; // 192
storage[798] =  11'b00011001010; // 202
storage[799] =  11'b00000001010; // 10
storage[800] =  11'b00011101101; // 237
storage[801] =  11'b00010100011; // 163
storage[802] = -11'b00010000000; // -128
storage[803] =  11'b00010110100; // 180
storage[804] =  11'b00010000011; // 131
storage[805] = -11'b00000010101; // -21
storage[806] =  11'b00011111011; // 251
storage[807] = -11'b00000000111; // -7
storage[808] = -11'b00000110011; // -51
storage[809] = -11'b00011000011; // -195
storage[810] = -11'b00000101010; // -42
storage[811] = -11'b00000111101; // -61
storage[812] =  11'b00011101100; // 236
storage[813] = -11'b00001001110; // -78
storage[814] = -11'b00001001001; // -73
storage[815] = -11'b00010000111; // -135
storage[816] =  11'b00001001000; // 72
storage[817] =  11'b00001010101; // 85
storage[818] = -11'b00000100010; // -34
storage[819] =  11'b00000010011; // 19
storage[820] =  11'b00011011101; // 221
storage[821] = -11'b00001000110; // -70
storage[822] = -11'b00001011101; // -93
storage[823] =  11'b00001100000; // 96
storage[824] = -11'b00011001011; // -203
storage[825] = -11'b00100001101; // -269
storage[826] = -11'b00000000110; // -6
storage[827] =  11'b00010101100; // 172
storage[828] = -11'b00011100011; // -227
storage[829] = -11'b00001110111; // -119
storage[830] = -11'b00001010111; // -87
storage[831] = -11'b00001001010; // -74
storage[832] = -11'b00011110011; // -243
storage[833] =  11'b00010101010; // 170
storage[834] = -11'b00000001110; // -14
storage[835] =  11'b00100001111; // 271
storage[836] =  11'b00011011100; // 220
storage[837] =  11'b00100101000; // 296
storage[838] = -11'b00001101001; // -105
storage[839] = -11'b00010111000; // -184
storage[840] = -11'b00000110010; // -50
storage[841] = -11'b00101001100; // -332
storage[842] = -11'b00011010101; // -213
storage[843] = -11'b00100011000; // -280
storage[844] = -11'b00001110111; // -119
storage[845] =  11'b00001011101; // 93
storage[846] = -11'b00000111000; // -56
storage[847] = -11'b00001000010; // -66
storage[848] =  11'b00000110010; // 50
storage[849] =  11'b00010001001; // 137
storage[850] = -11'b00101100010; // -354
storage[851] = -11'b01000010010; // -530
storage[852] = -11'b00011011000; // -216
storage[853] = -11'b00011011100; // -220
storage[854] = -11'b01101101010; // -874
storage[855] = -11'b00101101101; // -365
storage[856] = -11'b00001001110; // -78
storage[857] = -11'b00010000111; // -135
storage[858] = -11'b00100010001; // -273
storage[859] = -11'b00100100101; // -293
storage[860] =  11'b00010100001; // 161
storage[861] =  11'b00010011111; // 159
storage[862] = -11'b00001101100; // -108
storage[863] =  11'b00011001101; // 205
storage[864] = -11'b00010011011; // -155
storage[865] =  11'b00011111101; // 253
storage[866] =  11'b00011101110; // 238
storage[867] =  11'b00000110101; // 53
storage[868] = -11'b00000110110; // -54
storage[869] =  11'b00001001100; // 76
storage[870] =  11'b00000111001; // 57
storage[871] =  11'b00011000111; // 199
storage[872] = -11'b00001000100; // -68
storage[873] = -11'b00100110111; // -311
storage[874] =  11'b00000010111; // 23
storage[875] = -11'b00000111100; // -60
storage[876] =  11'b00000000100; // 4
storage[877] =  11'b00100111000; // 312
storage[878] =  11'b00011110110; // 246
storage[879] = -11'b00010011011; // -155
storage[880] =  11'b00000110111; // 55
storage[881] = -11'b00110011111; // -415
storage[882] =  11'b00001011000; // 88
storage[883] =  11'b00111101110; // 494
storage[884] =  11'b00000110010; // 50
storage[885] = -11'b00100110101; // -309
storage[886] = -11'b00001110110; // -118
storage[887] =  11'b00001001101; // 77
storage[888] =  11'b00100100010; // 290
storage[889] = -11'b00001111100; // -124
storage[890] = -11'b00001100110; // -102
storage[891] = -11'b00001010100; // -84
storage[892] = -11'b00010100001; // -161
storage[893] =  11'b00011010011; // 211
storage[894] =  11'b00010101000; // 168
storage[895] =  11'b00011110011; // 243
storage[896] =  11'b00001010000; // 80
storage[897] =  11'b00101001010; // 330
storage[898] =  11'b00011011111; // 223
storage[899] =  11'b00010010010; // 146
storage[900] =  11'b00011001111; // 207
storage[901] =  11'b00010011110; // 158
storage[902] =  11'b00001000101; // 69
storage[903] = -11'b00001100000; // -96
storage[904] =  11'b00010010010; // 146
storage[905] = -11'b00010000111; // -135
storage[906] = -11'b00000000100; // -4
storage[907] = -11'b00000011010; // -26
storage[908] = -11'b00001111101; // -125
storage[909] = -11'b00000101100; // -44
storage[910] = -11'b00001100101; // -101
storage[911] = -11'b00000001100; // -12
storage[912] = -11'b00101001001; // -329
storage[913] = -11'b00000010000; // -16
storage[914] =  11'b00010000101; // 133
storage[915] = -11'b00110101100; // -428
storage[916] =  11'b00001100101; // 101
storage[917] =  11'b00001010011; // 83
storage[918] = -11'b00111001101; // -461
storage[919] =  11'b00010010100; // 148
storage[920] =  11'b00011100011; // 227
storage[921] =  11'b00000011101; // 29
storage[922] =  11'b00011010101; // 213
storage[923] = -11'b00011101111; // -239
storage[924] = -11'b01010111100; // -700
storage[925] =  11'b00000110000; // 48
storage[926] =  11'b00000010000; // 16
storage[927] = -11'b00111101101; // -493
storage[928] = -11'b00011001010; // -202
storage[929] =  11'b00001000001; // 65
storage[930] =  11'b00011011100; // 220
storage[931] = -11'b00111110010; // -498
storage[932] = -11'b00101111100; // -380
storage[933] =  11'b00010100011; // 163
storage[934] = -11'b01001110100; // -628
storage[935] = -11'b00011101001; // -233
storage[936] = -11'b00000011111; // -31
storage[937] =  11'b00010001110; // 142
storage[938] = -11'b00010000110; // -134
storage[939] = -11'b00000010011; // -19
storage[940] =  11'b00010101101; // 173
storage[941] = -11'b00000110111; // -55
storage[942] =  11'b00011001100; // 204
storage[943] = -11'b00100011011; // -283
storage[944] = -11'b00010110111; // -183
storage[945] = -11'b00010110111; // -183
storage[946] =  11'b00010111110; // 190
storage[947] =  11'b00101100110; // 358
storage[948] =  11'b00001110011; // 115
storage[949] =  11'b00100010010; // 274
storage[950] =  11'b00110101110; // 430
storage[951] =  11'b00110011111; // 415
storage[952] =  11'b00001111000; // 120
storage[953] =  11'b00011100111; // 231
storage[954] =  11'b00001110101; // 117
storage[955] = -11'b00001010100; // -84
storage[956] = -11'b00110001010; // -394
storage[957] = -11'b00011001011; // -203
storage[958] =  11'b00111110001; // 497
storage[959] = -11'b00010110011; // -179
storage[960] =  11'b00001000100; // 68
storage[961] =  11'b00001001101; // 77
storage[962] =  11'b00100011101; // 285
storage[963] = -11'b00010100111; // -167
storage[964] =  11'b00000111001; // 57
storage[965] = -11'b00001010000; // -80
storage[966] =  11'b00000000110; // 6
storage[967] =  11'b00100011000; // 280
storage[968] =  11'b00101011000; // 344
storage[969] =  11'b00101011001; // 345
storage[970] =  11'b00010110001; // 177
storage[971] =  11'b00110100100; // 420
storage[972] =  11'b00010001011; // 139
storage[973] =  11'b00001010101; // 85
storage[974] =  11'b00001001011; // 75
storage[975] = -11'b00001110010; // -114
storage[976] = -11'b00010110110; // -182
storage[977] = -11'b00001001001; // -73
storage[978] = -11'b00010000011; // -131
storage[979] = -11'b00010010001; // -145
storage[980] =  11'b00001001010; // 74
storage[981] =  11'b00000000100; // 4
storage[982] = -11'b00000101010; // -42
storage[983] =  11'b00010000000; // 128
storage[984] =  11'b00011011111; // 223
storage[985] =  11'b00000100000; // 32
storage[986] =  11'b00011111101; // 253
storage[987] = -11'b00001100001; // -97
storage[988] =  11'b00011001011; // 203
storage[989] = -11'b00000010110; // -22
storage[990] = -11'b00011011101; // -221
storage[991] =  11'b00001101110; // 110
storage[992] =  11'b00000010000; // 16
storage[993] =  11'b00000001010; // 10
storage[994] =  11'b00000010111; // 23
storage[995] =  11'b00000111011; // 59
storage[996] =  11'b00001001011; // 75
storage[997] = -11'b00010110010; // -178
storage[998] = -11'b00010110111; // -183
storage[999] =  11'b00001100100; // 100
storage[1000] =  11'b00000101111; // 47
storage[1001] =  11'b00010001111; // 143
storage[1002] =  11'b00001110111; // 119
storage[1003] =  11'b00010001100; // 140
storage[1004] = -11'b00000001011; // -11
storage[1005] =  11'b00000111001; // 57
storage[1006] = -11'b00011100110; // -230
storage[1007] = -11'b00100111110; // -318
storage[1008] = -11'b00100010101; // -277
storage[1009] =  11'b00001001110; // 78
storage[1010] =  11'b00000101101; // 45
storage[1011] =  11'b00000010111; // 23
storage[1012] =  11'b00000111011; // 59
storage[1013] =  11'b00010001101; // 141
storage[1014] =  11'b00001110010; // 114
storage[1015] =  11'b00000101000; // 40
storage[1016] = -11'b00000001100; // -12
storage[1017] = -11'b00000100011; // -35
storage[1018] =  11'b00000011011; // 27
storage[1019] = -11'b00001101011; // -107
storage[1020] = -11'b00010011011; // -155
storage[1021] =  11'b00101011011; // 347
storage[1022] =  11'b00011010110; // 214
storage[1023] =  11'b00010110110; // 182
storage[1024] =  11'b00011111111; // 255
storage[1025] =  11'b00101100110; // 358
storage[1026] =  11'b00011100101; // 229
storage[1027] =  11'b00001000001; // 65
storage[1028] =  11'b00011011000; // 216
storage[1029] =  11'b00011001001; // 201
storage[1030] = -11'b00010001010; // -138
storage[1031] = -11'b00000101010; // -42
storage[1032] =  11'b00000100110; // 38
storage[1033] =  11'b00000101110; // 46
storage[1034] = -11'b00001100111; // -103
storage[1035] = -11'b00000100100; // -36
storage[1036] = -11'b00001001010; // -74
storage[1037] = -11'b00001010011; // -83
storage[1038] =  11'b00011011101; // 221
storage[1039] = -11'b00000011110; // -30
storage[1040] =  11'b00011010111; // 215
storage[1041] =  11'b00011101101; // 237
storage[1042] = -11'b00000110011; // -51
storage[1043] =  11'b00011111000; // 248
storage[1044] = -11'b00000110001; // -49
storage[1045] = -11'b00101101000; // -360
storage[1046] = -11'b00011110001; // -241
storage[1047] =  11'b00011110111; // 247
storage[1048] =  11'b00000010111; // 23
storage[1049] = -11'b00010001001; // -137
storage[1050] =  11'b00100010000; // 272
storage[1051] = -11'b00000001100; // -12
storage[1052] =  11'b00000111000; // 56
storage[1053] =  11'b00010000111; // 135
storage[1054] = -11'b00000010101; // -21
storage[1055] = -11'b00100001110; // -270
storage[1056] =  11'b00010101111; // 175
storage[1057] =  11'b00001110111; // 119
storage[1058] = -11'b00111010100; // -468
storage[1059] = -11'b00101100011; // -355
storage[1060] =  11'b00000010000; // 16
storage[1061] = -11'b00101101100; // -364
storage[1062] = -11'b00110001100; // -396
storage[1063] = -11'b00000011001; // -25
storage[1064] =  11'b00000010011; // 19
storage[1065] =  11'b00000111000; // 56
storage[1066] =  11'b00000101000; // 40
storage[1067] =  11'b00001010111; // 87
storage[1068] =  11'b00011100101; // 229
storage[1069] =  11'b00010001000; // 136
storage[1070] =  11'b00010010110; // 150
storage[1071] =  11'b00111011000; // 472
storage[1072] = -11'b00001111000; // -120
storage[1073] =  11'b00010000110; // 134
storage[1074] =  11'b00010011001; // 153
storage[1075] = -11'b00100011101; // -285
storage[1076] = -11'b00011001111; // -207
storage[1077] = -11'b00001001110; // -78
storage[1078] = -11'b00001100100; // -100
storage[1079] =  11'b00010110101; // 181
storage[1080] =  11'b00011001101; // 205
storage[1081] = -11'b00000101101; // -45
storage[1082] =  11'b00011110100; // 244
storage[1083] =  11'b00010010011; // 147
storage[1084] = -11'b00000011111; // -31
storage[1085] = -11'b00000110001; // -49
storage[1086] = -11'b00000010111; // -23
storage[1087] = -11'b00010010001; // -145
storage[1088] = -11'b00000101100; // -44
storage[1089] = -11'b00011101000; // -232
storage[1090] = -11'b00010101100; // -172
storage[1091] = -11'b00100000001; // -257
storage[1092] = -11'b00000110001; // -49
storage[1093] = -11'b00001010010; // -82
storage[1094] = -11'b00011011110; // -222
storage[1095] =  11'b00001100110; // 102
storage[1096] =  11'b00100000110; // 262
storage[1097] =  11'b00011101000; // 232
storage[1098] = -11'b00000001001; // -9
storage[1099] =  11'b00000110100; // 52
storage[1100] =  11'b00001110011; // 115
storage[1101] = -11'b00010001111; // -143
storage[1102] =  11'b00100101111; // 303
storage[1103] =  11'b00100010001; // 273
storage[1104] =  11'b00000010101; // 21
storage[1105] =  11'b00000101110; // 46
storage[1106] =  11'b00101001111; // 335
storage[1107] =  11'b00000011001; // 25
storage[1108] =  11'b00000110010; // 50
storage[1109] =  11'b00010011000; // 152
storage[1110] = -11'b00000111000; // -56
storage[1111] = -11'b00010100001; // -161
storage[1112] = -11'b00010001100; // -140
storage[1113] =  11'b00011011101; // 221
storage[1114] =  11'b00010000001; // 129
storage[1115] = -11'b00001110101; // -117
storage[1116] =  11'b00011011100; // 220
storage[1117] = -11'b00000111110; // -62
storage[1118] =  11'b00001001101; // 77
storage[1119] = -11'b00001000100; // -68
storage[1120] = -11'b00001110100; // -116
storage[1121] =  11'b00000010100; // 20
storage[1122] =  11'b00000100000; // 32
storage[1123] =  11'b00000000010; // 2
storage[1124] = -11'b00010011010; // -154
storage[1125] =  11'b00001011111; // 95
storage[1126] = -11'b00101011110; // -350
storage[1127] =  11'b00000010000; // 16
storage[1128] =  11'b00001111100; // 124
storage[1129] =  11'b00001011001; // 89
storage[1130] =  11'b00101010011; // 339
storage[1131] =  11'b00100010000; // 272
storage[1132] = -11'b00000101001; // -41
storage[1133] =  11'b00011000001; // 193
storage[1134] =  11'b00100011001; // 281
storage[1135] = -11'b00010001000; // -136
storage[1136] = -11'b00001011101; // -93
storage[1137] =  11'b00000010001; // 17
storage[1138] =  11'b00000111101; // 61
storage[1139] = -11'b00000011111; // -31
storage[1140] = -11'b00001100011; // -99
storage[1141] =  11'b00001010011; // 83
storage[1142] = -11'b00000000011; // -3
storage[1143] =  11'b00000010000; // 16
storage[1144] = -11'b00011001101; // -205
storage[1145] = -11'b00010101100; // -172
storage[1146] = -11'b00000100100; // -36
storage[1147] = -11'b00010111101; // -189
storage[1148] = -11'b00111001010; // -458
storage[1149] = -11'b00000001101; // -13
storage[1150] = -11'b00011011010; // -218
storage[1151] = -11'b00010110100; // -180
storage[1152] = -11'b00000000111; // -7
storage[1153] =  11'b00001010001; // 81
storage[1154] =  11'b00011001011; // 203
storage[1155] = -11'b00000010110; // -22
storage[1156] =  11'b00011110100; // 244
storage[1157] =  11'b00101010011; // 339
storage[1158] =  11'b00001001100; // 76
storage[1159] = -11'b00000001101; // -13
storage[1160] =  11'b00000101110; // 46
storage[1161] =  11'b00000011110; // 30
storage[1162] = -11'b00011011011; // -219
storage[1163] =  11'b00000000011; // 3
storage[1164] =  11'b00011010000; // 208
storage[1165] = -11'b01001011010; // -602
storage[1166] = -11'b00000101101; // -45
storage[1167] =  11'b00010101011; // 171
storage[1168] = -11'b00011111110; // -254
storage[1169] =  11'b00011110101; // 245
storage[1170] =  11'b00011010010; // 210
storage[1171] = -11'b00100010100; // -276
storage[1172] = -11'b00010111111; // -191
storage[1173] = -11'b00100011011; // -283
storage[1174] = -11'b00000010110; // -22
storage[1175] =  11'b00000010011; // 19
storage[1176] =  11'b00000011110; // 30
storage[1177] =  11'b00100011111; // 287
storage[1178] =  11'b00000100111; // 39
storage[1179] = -11'b00001001111; // -79
storage[1180] =  11'b00001000010; // 66
storage[1181] = -11'b00000010001; // -17
storage[1182] =  11'b00001001111; // 79
storage[1183] =  11'b00001111011; // 123
storage[1184] =  11'b00001100011; // 99
storage[1185] = -11'b00010100111; // -167
storage[1186] = -11'b00001011110; // -94
storage[1187] = -11'b00000100111; // -39
storage[1188] = -11'b00101000011; // -323
storage[1189] =  11'b00000111001; // 57
storage[1190] = -11'b00000100000; // -32
storage[1191] =  11'b00010010001; // 145
storage[1192] =  11'b00001010100; // 84
storage[1193] = -11'b00010100010; // -162
storage[1194] = -11'b00001010001; // -81
storage[1195] =  11'b00001011000; // 88
storage[1196] = -11'b00001010101; // -85
storage[1197] = -11'b00010111000; // -184
storage[1198] = -11'b00001011001; // -89
storage[1199] = -11'b00001000011; // -67
storage[1200] =  11'b00011101110; // 238
storage[1201] =  11'b00001110111; // 119
storage[1202] =  11'b00000110101; // 53
storage[1203] =  11'b00100001010; // 266
storage[1204] = -11'b00000101011; // -43
storage[1205] =  11'b00001011111; // 95
storage[1206] =  11'b00100011110; // 286
storage[1207] = -11'b00001011011; // -91
storage[1208] =  11'b00100110000; // 304
storage[1209] = -11'b00010100001; // -161
storage[1210] =  11'b00000011111; // 31
storage[1211] =  11'b00011000101; // 197
storage[1212] = -11'b00001001100; // -76
storage[1213] = -11'b00000111111; // -63
storage[1214] = -11'b00000011000; // -24
storage[1215] = -11'b00010100110; // -166
storage[1216] = -11'b00001010001; // -81
storage[1217] =  11'b00010010011; // 147
storage[1218] =  11'b00100001010; // 266
storage[1219] =  11'b00001010101; // 85
storage[1220] = -11'b00000100001; // -33
storage[1221] = -11'b00001100000; // -96
storage[1222] = -11'b00001000001; // -65
storage[1223] = -11'b00001000101; // -69
storage[1224] = -11'b00001110010; // -114
storage[1225] = -11'b00000110001; // -49
storage[1226] =  11'b00000000001; // 1
storage[1227] = -11'b00000101111; // -47
storage[1228] = -11'b00000110111; // -55
storage[1229] = -11'b00001000010; // -66
storage[1230] = -11'b00000111110; // -62
storage[1231] =  11'b00000010100; // 20
storage[1232] = -11'b00011101110; // -238
storage[1233] =  11'b00000000111; // 7
storage[1234] = -11'b00000110101; // -53
storage[1235] =  11'b00101110101; // 373
storage[1236] =  11'b00011011001; // 217
storage[1237] =  11'b00000111101; // 61
storage[1238] = -11'b00000010101; // -21
storage[1239] = -11'b00001101111; // -111
storage[1240] = -11'b00010010010; // -146
storage[1241] = -11'b00001100101; // -101
storage[1242] = -11'b00001110000; // -112
storage[1243] =  11'b00001110101; // 117
storage[1244] =  11'b00111001000; // 456
storage[1245] =  11'b00010011111; // 159
storage[1246] = -11'b00000101010; // -42
storage[1247] = -11'b00001111000; // -120
storage[1248] =  11'b00010110010; // 178
storage[1249] =  11'b00000000101; // 5
storage[1250] = -11'b00010110011; // -179
storage[1251] =  11'b00001011000; // 88
storage[1252] = -11'b00100001111; // -271
storage[1253] = -11'b00100000001; // -257
storage[1254] = -11'b00011011011; // -219
storage[1255] =  11'b00010001100; // 140
storage[1256] =  11'b00000100100; // 36
storage[1257] =  11'b00010000100; // 132
storage[1258] =  11'b00000110111; // 55
storage[1259] = -11'b00000000010; // -2
storage[1260] =  11'b00001111011; // 123
storage[1261] =  11'b00000010011; // 19
storage[1262] =  11'b00001000110; // 70
storage[1263] =  11'b00001010100; // 84
storage[1264] = -11'b00010100100; // -164
storage[1265] = -11'b00010110111; // -183
storage[1266] = -11'b00000110110; // -54
storage[1267] =  11'b00010110101; // 181
storage[1268] =  11'b00001010101; // 85
storage[1269] =  11'b00010101100; // 172
storage[1270] = -11'b00000010111; // -23
storage[1271] = -11'b00000011110; // -30
storage[1272] = -11'b00000001011; // -11
storage[1273] =  11'b00000001111; // 15
storage[1274] = -11'b00001010000; // -80
storage[1275] =  11'b00000111000; // 56
storage[1276] =  11'b00001000011; // 67
storage[1277] = -11'b00001010110; // -86
storage[1278] = -11'b00000011000; // -24
storage[1279] =  11'b00000000010; // 2
storage[1280] = -11'b00001010011; // -83
storage[1281] = -11'b00001001010; // -74
storage[1282] =  11'b00011000100; // 196
storage[1283] =  11'b00001111011; // 123
storage[1284] =  11'b00001011001; // 89
storage[1285] =  11'b00000011100; // 28
storage[1286] = -11'b00001110101; // -117
storage[1287] = -11'b00001001100; // -76
storage[1288] = -11'b00010011010; // -154
storage[1289] = -11'b00010000100; // -132
storage[1290] = -11'b00001100110; // -102
storage[1291] = -11'b00011110111; // -247
storage[1292] = -11'b00010100110; // -166
storage[1293] = -11'b00001010011; // -83
storage[1294] = -11'b00010110100; // -180
storage[1295] = -11'b00010001000; // -136
storage[1296] = -11'b00001110000; // -112
storage[1297] =  11'b00000111100; // 60
storage[1298] = -11'b00000011101; // -29
storage[1299] = -11'b00001010110; // -86
storage[1300] =  11'b00000001000; // 8
storage[1301] = -11'b00001011111; // -95
storage[1302] = -11'b00000010010; // -18
storage[1303] = -11'b00010100111; // -167
storage[1304] = -11'b00100000001; // -257
storage[1305] = -11'b00010110010; // -178
storage[1306] =  11'b00010001110; // 142
storage[1307] =  11'b00011100001; // 225
storage[1308] = -11'b00001100011; // -99
storage[1309] =  11'b00000100111; // 39
storage[1310] =  11'b00000100101; // 37
storage[1311] = -11'b00011100101; // -229
storage[1312] =  11'b00001101111; // 111
storage[1313] =  11'b00001010100; // 84
storage[1314] =  11'b00001010111; // 87
storage[1315] =  11'b00000100101; // 37
storage[1316] =  11'b00001011010; // 90
storage[1317] =  11'b00011001111; // 207
storage[1318] =  11'b00001010101; // 85
storage[1319] =  11'b00001001100; // 76
storage[1320] =  11'b00011010101; // 213
storage[1321] =  11'b00000101000; // 40
storage[1322] =  11'b00000010000; // 16
storage[1323] =  11'b00001011000; // 88
storage[1324] =  11'b00000000000; // 0
storage[1325] = -11'b00000010101; // -21
storage[1326] = -11'b00010111101; // -189
storage[1327] = -11'b00001011010; // -90
storage[1328] =  11'b00000011010; // 26
storage[1329] = -11'b00001100100; // -100
storage[1330] =  11'b00010000011; // 131
storage[1331] =  11'b00001100010; // 98
storage[1332] = -11'b00001011110; // -94
storage[1333] = -11'b00001011100; // -92
storage[1334] = -11'b00000010110; // -22
storage[1335] = -11'b00000001001; // -9
storage[1336] = -11'b00000000010; // -2
storage[1337] = -11'b00000010100; // -20
storage[1338] =  11'b00000010010; // 18
storage[1339] =  11'b00001100111; // 103
storage[1340] =  11'b00000011101; // 29
storage[1341] =  11'b00000010001; // 17
storage[1342] = -11'b00000110100; // -52
storage[1343] =  11'b00000010000; // 16
storage[1344] = -11'b00000100101; // -37
storage[1345] = -11'b00000010000; // -16
storage[1346] =  11'b00001110101; // 117
storage[1347] =  11'b00000110001; // 49
storage[1348] =  11'b00010011001; // 153
storage[1349] =  11'b00010010111; // 151
storage[1350] =  11'b00000011101; // 29
storage[1351] = -11'b00000111001; // -57
storage[1352] =  11'b00000000011; // 3
storage[1353] =  11'b00000010101; // 21
storage[1354] = -11'b00001001100; // -76
storage[1355] =  11'b00000000111; // 7
storage[1356] = -11'b00001011010; // -90
storage[1357] = -11'b00000011001; // -25
storage[1358] = -11'b00001011110; // -94
storage[1359] = -11'b00000111010; // -58
storage[1360] =  11'b00001100010; // 98
storage[1361] =  11'b00010001000; // 136
storage[1362] =  11'b00001011111; // 95
storage[1363] =  11'b00010010101; // 149
storage[1364] =  11'b00100001010; // 266
storage[1365] =  11'b00001010101; // 85
storage[1366] =  11'b00001110000; // 112
storage[1367] = -11'b00000110111; // -55
storage[1368] = -11'b00000111000; // -56
storage[1369] = -11'b00000101010; // -42
storage[1370] = -11'b00001000010; // -66
storage[1371] = -11'b00000001011; // -11
storage[1372] =  11'b00001010111; // 87
storage[1373] = -11'b00000011100; // -28
storage[1374] =  11'b00000000101; // 5
storage[1375] = -11'b00000000111; // -7
storage[1376] =  11'b00000100000; // 32
storage[1377] =  11'b00001000111; // 71
storage[1378] = -11'b00001011100; // -92
storage[1379] = -11'b00001000001; // -65
storage[1380] = -11'b00000111000; // -56
storage[1381] = -11'b00001101111; // -111
storage[1382] =  11'b00000101001; // 41
storage[1383] = -11'b00001110100; // -116
storage[1384] =  11'b00001100100; // 100
storage[1385] = -11'b00000000110; // -6
storage[1386] =  11'b00000011100; // 28
storage[1387] =  11'b00000101100; // 44
storage[1388] =  11'b00001111011; // 123
storage[1389] =  11'b00001011100; // 92
storage[1390] =  11'b00010100111; // 167
storage[1391] =  11'b00011111010; // 250
storage[1392] =  11'b00000000100; // 4
storage[1393] =  11'b00011111000; // 248
storage[1394] =  11'b00011110110; // 246
storage[1395] =  11'b00100000100; // 260
storage[1396] = -11'b00011100110; // -230
storage[1397] =  11'b00000010011; // 19
storage[1398] =  11'b00000000111; // 7
storage[1399] = -11'b00000100110; // -38
storage[1400] =  11'b00000000010; // 2
storage[1401] =  11'b00000000010; // 2
storage[1402] = -11'b00001000011; // -67
storage[1403] =  11'b00001011111; // 95
storage[1404] =  11'b00001010110; // 86
storage[1405] = -11'b00000111010; // -58
storage[1406] = -11'b00000010001; // -17
storage[1407] = -11'b00001111000; // -120
storage[1408] =  11'b00001100010; // 98
storage[1409] = -11'b00000101100; // -44
storage[1410] = -11'b00010011111; // -159
storage[1411] =  11'b00010110001; // 177
storage[1412] =  11'b00000110100; // 52
storage[1413] = -11'b00000011010; // -26
storage[1414] =  11'b00001000110; // 70
storage[1415] = -11'b00001100011; // -99
storage[1416] = -11'b00000010010; // -18
storage[1417] =  11'b00010011001; // 153
storage[1418] = -11'b00000110100; // -52
storage[1419] = -11'b00000011110; // -30
storage[1420] =  11'b00001100111; // 103
storage[1421] =  11'b00001011001; // 89
storage[1422] =  11'b00000010111; // 23
storage[1423] =  11'b00001010110; // 86
storage[1424] = -11'b00000011101; // -29
storage[1425] = -11'b00010110011; // -179
storage[1426] =  11'b00000011101; // 29
storage[1427] =  11'b00001101100; // 108
storage[1428] =  11'b00001000100; // 68
storage[1429] = -11'b00001110110; // -118
storage[1430] =  11'b00001101100; // 108
storage[1431] =  11'b00011110100; // 244
storage[1432] = -11'b00011110011; // -243
storage[1433] = -11'b00000000100; // -4
storage[1434] = -11'b00000010111; // -23
storage[1435] = -11'b00011100001; // -225
storage[1436] = -11'b00001100101; // -101
storage[1437] =  11'b00001101010; // 106
storage[1438] =  11'b00011111000; // 248
storage[1439] = -11'b00101010100; // -340
storage[1440] =  11'b00000110111; // 55
storage[1441] = -11'b00001111111; // -127
storage[1442] =  11'b00000010000; // 16
storage[1443] =  11'b00001111000; // 120
storage[1444] = -11'b00100011001; // -281
storage[1445] = -11'b00010001001; // -137
storage[1446] =  11'b00010000001; // 129
storage[1447] = -11'b00001000111; // -71
storage[1448] = -11'b00111000000; // -448
storage[1449] =  11'b00000000011; // 3
storage[1450] =  11'b00000110110; // 54
storage[1451] = -11'b00000000101; // -5
storage[1452] = -11'b00001110111; // -119
storage[1453] =  11'b00001011011; // 91
storage[1454] =  11'b00001000000; // 64
storage[1455] = -11'b00010000110; // -134
storage[1456] =  11'b00001110010; // 114
storage[1457] =  11'b00010101100; // 172
storage[1458] =  11'b00000000010; // 2
storage[1459] =  11'b00010110111; // 183
storage[1460] =  11'b00001010101; // 85
storage[1461] =  11'b00010010001; // 145
storage[1462] =  11'b00101001010; // 330
storage[1463] =  11'b00000011100; // 28
storage[1464] =  11'b00001100010; // 98
storage[1465] =  11'b00010100100; // 164
storage[1466] =  11'b00001010001; // 81
storage[1467] = -11'b00000100011; // -35
storage[1468] = -11'b00000101011; // -43
storage[1469] =  11'b00000110101; // 53
storage[1470] =  11'b00010101010; // 170
storage[1471] = -11'b00001101101; // -109
storage[1472] =  11'b00000000110; // 6
storage[1473] =  11'b00001001010; // 74
storage[1474] = -11'b00000110000; // -48
storage[1475] = -11'b00000011001; // -25
storage[1476] =  11'b00000101101; // 45
storage[1477] =  11'b00000000110; // 6
storage[1478] = -11'b00001011011; // -91
storage[1479] =  11'b00000001000; // 8
storage[1480] =  11'b00000011110; // 30
storage[1481] =  11'b00000100100; // 36
storage[1482] =  11'b00010011101; // 157
storage[1483] = -11'b00000110011; // -51
storage[1484] = -11'b00000110111; // -55
storage[1485] =  11'b00010000011; // 131
storage[1486] =  11'b00001101110; // 110
storage[1487] =  11'b00001100001; // 97
storage[1488] =  11'b00001111110; // 126
storage[1489] =  11'b00000000011; // 3
storage[1490] =  11'b00001010110; // 86
storage[1491] = -11'b00001110111; // -119
storage[1492] = -11'b00000101111; // -47
storage[1493] =  11'b00000011000; // 24
storage[1494] = -11'b00000110000; // -48
storage[1495] =  11'b00001100000; // 96
storage[1496] =  11'b00011001001; // 201
storage[1497] =  11'b00001010010; // 82
storage[1498] = -11'b00000101000; // -40
storage[1499] = -11'b00000000100; // -4
storage[1500] =  11'b00000110110; // 54
storage[1501] = -11'b00000011001; // -25
storage[1502] = -11'b00001111101; // -125
storage[1503] =  11'b00000110010; // 50
storage[1504] = -11'b00011011011; // -219
storage[1505] =  11'b00000111011; // 59
storage[1506] = -11'b00000001110; // -14
storage[1507] = -11'b00000000100; // -4
storage[1508] = -11'b00000110000; // -48
storage[1509] =  11'b00001010111; // 87
storage[1510] =  11'b00001100101; // 101
storage[1511] =  11'b00011101000; // 232
storage[1512] =  11'b00011101010; // 234
storage[1513] = -11'b00010101011; // -171
storage[1514] = -11'b00011010100; // -212
storage[1515] = -11'b00010110110; // -182
storage[1516] =  11'b00000011010; // 26
storage[1517] = -11'b00101101000; // -360
storage[1518] = -11'b00010010011; // -147
storage[1519] =  11'b00001100110; // 102
storage[1520] =  11'b00000011001; // 25
storage[1521] = -11'b00001010111; // -87
storage[1522] = -11'b00001100000; // -96
storage[1523] =  11'b00011100111; // 231
storage[1524] =  11'b00000110100; // 52
storage[1525] = -11'b00010110101; // -181
storage[1526] =  11'b00001001000; // 72
storage[1527] =  11'b00010111000; // 184
storage[1528] = -11'b00000110011; // -51
storage[1529] = -11'b00011101001; // -233
storage[1530] = -11'b00000100111; // -39
storage[1531] = -11'b00001001110; // -78
storage[1532] =  11'b00001010010; // 82
storage[1533] =  11'b00001101011; // 107
storage[1534] = -11'b00000100000; // -32
storage[1535] =  11'b00010001101; // 141
storage[1536] =  11'b00010000011; // 131
storage[1537] = -11'b00000110110; // -54
storage[1538] =  11'b00000011110; // 30
storage[1539] = -11'b00010000101; // -133
storage[1540] = -11'b00001100111; // -103
storage[1541] = -11'b00011001001; // -201
storage[1542] = -11'b00001111001; // -121
storage[1543] = -11'b00000011000; // -24
storage[1544] = -11'b00001011101; // -93
storage[1545] =  11'b00000000010; // 2
storage[1546] =  11'b00000100110; // 38
storage[1547] =  11'b00000010110; // 22
storage[1548] = -11'b00000100000; // -32
storage[1549] =  11'b00000010110; // 22
storage[1550] = -11'b00000110100; // -52
storage[1551] =  11'b00000010000; // 16
storage[1552] =  11'b00010010110; // 150
storage[1553] = -11'b00000101111; // -47
storage[1554] = -11'b00000101001; // -41
storage[1555] =  11'b00001111110; // 126
storage[1556] =  11'b00000010001; // 17
storage[1557] = -11'b00001001010; // -74
storage[1558] =  11'b00000010101; // 21
storage[1559] = -11'b00000000010; // -2
storage[1560] =  11'b00000101101; // 45
storage[1561] = -11'b00001100011; // -99
storage[1562] = -11'b00010001110; // -142
storage[1563] = -11'b00000100110; // -38
storage[1564] = -11'b00010000110; // -134
storage[1565] = -11'b00000110110; // -54
storage[1566] =  11'b00001010010; // 82
storage[1567] =  11'b00000010101; // 21
storage[1568] = -11'b00000011010; // -26
storage[1569] =  11'b00001100100; // 100
storage[1570] =  11'b00010001111; // 143
storage[1571] =  11'b00000011111; // 31
storage[1572] =  11'b00001110110; // 118
storage[1573] = -11'b00000101010; // -42
storage[1574] =  11'b00000001100; // 12
storage[1575] =  11'b00001111100; // 124
storage[1576] =  11'b00000000100; // 4
storage[1577] = -11'b00001000010; // -66
storage[1578] = -11'b00011011101; // -221
storage[1579] =  11'b00000001011; // 11
storage[1580] =  11'b00000001011; // 11
storage[1581] =  11'b00010010010; // 146
storage[1582] =  11'b00001011000; // 88
storage[1583] =  11'b00010110011; // 179
storage[1584] =  11'b00010010010; // 146
storage[1585] =  11'b00001010101; // 85
storage[1586] = -11'b00000001100; // -12
storage[1587] = -11'b00000111000; // -56
storage[1588] =  11'b00000011000; // 24
storage[1589] =  11'b00000110011; // 51
storage[1590] =  11'b00000100011; // 35
storage[1591] =  11'b00000110111; // 55
storage[1592] = -11'b00000001010; // -10
storage[1593] = -11'b00000011111; // -31
storage[1594] = -11'b00000100100; // -36
storage[1595] =  11'b00000101101; // 45
storage[1596] = -11'b00001010110; // -86
storage[1597] =  11'b00000010001; // 17
storage[1598] =  11'b00000011011; // 27
storage[1599] =  11'b00001001001; // 73
storage[1600] =  11'b00010011011; // 155
storage[1601] =  11'b00100011110; // 286
storage[1602] =  11'b00011000110; // 198
storage[1603] =  11'b00001111111; // 127
storage[1604] =  11'b00100010100; // 276
storage[1605] =  11'b00101001100; // 332
storage[1606] =  11'b00000111000; // 56
storage[1607] =  11'b00001100011; // 99
storage[1608] =  11'b00100110011; // 307
storage[1609] =  11'b00101010111; // 343
storage[1610] =  11'b00100111011; // 315
storage[1611] =  11'b00100101011; // 299
storage[1612] =  11'b00000001100; // 12
storage[1613] =  11'b00000111110; // 62
storage[1614] =  11'b00000000001; // 1
storage[1615] =  11'b00011000011; // 195
storage[1616] =  11'b00011101010; // 234
storage[1617] =  11'b00010010010; // 146
storage[1618] =  11'b00001101110; // 110
storage[1619] =  11'b00000010111; // 23
storage[1620] = -11'b00000110100; // -52
storage[1621] = -11'b00000000101; // -5
storage[1622] = -11'b00000110101; // -53
storage[1623] = -11'b00000111101; // -61
storage[1624] =  11'b00000011101; // 29
storage[1625] = -11'b00000100001; // -33
storage[1626] =  11'b00000110010; // 50
storage[1627] =  11'b00000011111; // 31
storage[1628] =  11'b00000110010; // 50
storage[1629] =  11'b00000101101; // 45
storage[1630] = -11'b00010011100; // -156
storage[1631] = -11'b00010100001; // -161
storage[1632] = -11'b00001101011; // -107
storage[1633] =  11'b00001110100; // 116
storage[1634] =  11'b00010001001; // 137
storage[1635] =  11'b00000010010; // 18
storage[1636] =  11'b00001101101; // 109
storage[1637] =  11'b00001000011; // 67
storage[1638] =  11'b00000001100; // 12
storage[1639] = -11'b00000001111; // -15
storage[1640] = -11'b00000100110; // -38
storage[1641] = -11'b00010001111; // -143
storage[1642] =  11'b00010010111; // 151
storage[1643] =  11'b00000001000; // 8
storage[1644] = -11'b00000001001; // -9
storage[1645] =  11'b00010101010; // 170
storage[1646] = -11'b00010101111; // -175
storage[1647] = -11'b00001100011; // -99
storage[1648] = -11'b00010010000; // -144
storage[1649] =  11'b00011100010; // 226
storage[1650] =  11'b00011001111; // 207
storage[1651] =  11'b00001000010; // 66
storage[1652] =  11'b00010000000; // 128
storage[1653] =  11'b00000111111; // 63
storage[1654] = -11'b00000010001; // -17
storage[1655] =  11'b00010001011; // 139
storage[1656] =  11'b00001001111; // 79
storage[1657] =  11'b00010001000; // 136
storage[1658] =  11'b00000000101; // 5
storage[1659] = -11'b00001000101; // -69
storage[1660] =  11'b00001001100; // 76
storage[1661] = -11'b00011110111; // -247
storage[1662] = -11'b00011011010; // -218
storage[1663] = -11'b00011100001; // -225
storage[1664] = -11'b00011111000; // -248
storage[1665] =  11'b00011000001; // 193
storage[1666] =  11'b00010100010; // 162
storage[1667] =  11'b00001010101; // 85
storage[1668] =  11'b00000010001; // 17
storage[1669] = -11'b00000110100; // -52
storage[1670] = -11'b00010101011; // -171
storage[1671] = -11'b00000111010; // -58
storage[1672] = -11'b00100010111; // -279
storage[1673] = -11'b00111100010; // -482
storage[1674] = -11'b00001100000; // -96
storage[1675] =  11'b00000001011; // 11
storage[1676] =  11'b00000111110; // 62
storage[1677] =  11'b00001100011; // 99
storage[1678] =  11'b00000100001; // 33
storage[1679] =  11'b00000100001; // 33
storage[1680] =  11'b00000010100; // 20
storage[1681] =  11'b00010010000; // 144
storage[1682] =  11'b00010001010; // 138
storage[1683] =  11'b00000001110; // 14
storage[1684] =  11'b00010100110; // 166
storage[1685] = -11'b00001011110; // -94
storage[1686] =  11'b00000010100; // 20
storage[1687] =  11'b00010111110; // 190
storage[1688] = -11'b00001010100; // -84
storage[1689] = -11'b00001010000; // -80
storage[1690] =  11'b00001100111; // 103
storage[1691] = -11'b00001010100; // -84
storage[1692] = -11'b00000110110; // -54
storage[1693] =  11'b00001001000; // 72
storage[1694] =  11'b00010000101; // 133
storage[1695] =  11'b00001000011; // 67
storage[1696] = -11'b00000111110; // -62
storage[1697] = -11'b00000101110; // -46
storage[1698] =  11'b00001001011; // 75
storage[1699] =  11'b00000010000; // 16
storage[1700] =  11'b00000111010; // 58
storage[1701] =  11'b00000100111; // 39
storage[1702] = -11'b00101101010; // -362
storage[1703] =  11'b00011010000; // 208
storage[1704] =  11'b00000011001; // 25
storage[1705] = -11'b00010000010; // -130
storage[1706] =  11'b00001001001; // 73
storage[1707] = -11'b00000100001; // -33
storage[1708] = -11'b00010001111; // -143
storage[1709] =  11'b00010110111; // 183
storage[1710] =  11'b00000011010; // 26
storage[1711] = -11'b00010010000; // -144
storage[1712] = -11'b00010010011; // -147
storage[1713] =  11'b00001100001; // 97
storage[1714] = -11'b00001111110; // -126
storage[1715] = -11'b00011101001; // -233
storage[1716] =  11'b00010110111; // 183
storage[1717] = -11'b00010101000; // -168
storage[1718] = -11'b00000111001; // -57
storage[1719] =  11'b00010111000; // 184
storage[1720] =  11'b00010011001; // 153
storage[1721] =  11'b00001111110; // 126
storage[1722] =  11'b00001110101; // 117
storage[1723] =  11'b00011000011; // 195
storage[1724] =  11'b00001100010; // 98
storage[1725] =  11'b00001100111; // 103
storage[1726] =  11'b00000011111; // 31
storage[1727] = -11'b00000011010; // -26
storage[1728] = -11'b00000111111; // -63
storage[1729] =  11'b00010110100; // 180
storage[1730] = -11'b00010101110; // -174
storage[1731] = -11'b00001101010; // -106
storage[1732] =  11'b00000110001; // 49
storage[1733] = -11'b00011000110; // -198
storage[1734] = -11'b00001110111; // -119
storage[1735] = -11'b00000000100; // -4
storage[1736] = -11'b00011010101; // -213
storage[1737] = -11'b00000110001; // -49
storage[1738] =  11'b00001001101; // 77
storage[1739] =  11'b00000111111; // 63
storage[1740] =  11'b00001010000; // 80
storage[1741] =  11'b00000011101; // 29
storage[1742] =  11'b00000101100; // 44
storage[1743] =  11'b00000000011; // 3
storage[1744] =  11'b00000000011; // 3
storage[1745] =  11'b00001000101; // 69
storage[1746] = -11'b00000010101; // -21
storage[1747] = -11'b00011111011; // -251
storage[1748] = -11'b00000000101; // -5
storage[1749] = -11'b00100000101; // -261
storage[1750] = -11'b00101010001; // -337
storage[1751] = -11'b00000110011; // -51
storage[1752] = -11'b00011001010; // -202
storage[1753] = -11'b00011011111; // -223
storage[1754] = -11'b00001011010; // -90
storage[1755] = -11'b00011100010; // -226
storage[1756] =  11'b00001000010; // 66
storage[1757] = -11'b00001010001; // -81
storage[1758] = -11'b00011001010; // -202
storage[1759] = -11'b00000111001; // -57
storage[1760] =  11'b00000100000; // 32
storage[1761] = -11'b00100000010; // -258
storage[1762] =  11'b00000100111; // 39
storage[1763] =  11'b00010001011; // 139
storage[1764] = -11'b00001110011; // -115
storage[1765] =  11'b00000010110; // 22
storage[1766] =  11'b00001001011; // 75
storage[1767] =  11'b00010010101; // 149
storage[1768] =  11'b00001010011; // 83
storage[1769] = -11'b00000111110; // -62
storage[1770] =  11'b00000101001; // 41
storage[1771] =  11'b00000110000; // 48
storage[1772] = -11'b00000111010; // -58
storage[1773] =  11'b00001010110; // 86
storage[1774] = -11'b00001110001; // -113
storage[1775] = -11'b00100101001; // -297
storage[1776] =  11'b00001001101; // 77
storage[1777] = -11'b00100100111; // -295
storage[1778] = -11'b00001110101; // -117
storage[1779] =  11'b00001101001; // 105
storage[1780] = -11'b00000101011; // -43
storage[1781] = -11'b00000011111; // -31
storage[1782] =  11'b00010101101; // 173
storage[1783] = -11'b00001011001; // -89
storage[1784] =  11'b00010101000; // 168
storage[1785] = -11'b00011010001; // -209
storage[1786] =  11'b00001100001; // 97
storage[1787] = -11'b00000110110; // -54
storage[1788] = -11'b00010100010; // -162
storage[1789] =  11'b00001100110; // 102
storage[1790] =  11'b00000000110; // 6
storage[1791] =  11'b00000101101; // 45
storage[1792] = -11'b00001100001; // -97
storage[1793] =  11'b00011011110; // 222
storage[1794] =  11'b00000110110; // 54
storage[1795] =  11'b00000100010; // 34
storage[1796] =  11'b00011111100; // 252
storage[1797] =  11'b00001111011; // 123
storage[1798] = -11'b00001011000; // -88
storage[1799] =  11'b00011001011; // 203
storage[1800] =  11'b00010011011; // 155
storage[1801] = -11'b00000111111; // -63
storage[1802] = -11'b00001010011; // -83
storage[1803] = -11'b00010111101; // -189
storage[1804] =  11'b00000011011; // 27
storage[1805] = -11'b00000011001; // -25
storage[1806] = -11'b00011110111; // -247
storage[1807] = -11'b00000000110; // -6
storage[1808] = -11'b00000010010; // -18
storage[1809] = -11'b00010011111; // -159
storage[1810] = -11'b00001011011; // -91
storage[1811] =  11'b00011011110; // 222
storage[1812] =  11'b00001010001; // 81
storage[1813] = -11'b00000100110; // -38
storage[1814] =  11'b00100001010; // 266
storage[1815] =  11'b00010000101; // 133
storage[1816] =  11'b00001101101; // 109
storage[1817] =  11'b00000111000; // 56
storage[1818] =  11'b00010000001; // 129
storage[1819] =  11'b00000010000; // 16
storage[1820] =  11'b00011000001; // 193
storage[1821] =  11'b00011011100; // 220
storage[1822] =  11'b00000000000; // 0
storage[1823] =  11'b00101111110; // 382
storage[1824] =  11'b00000101101; // 45
storage[1825] =  11'b00011110111; // 247
storage[1826] =  11'b00110000110; // 390
storage[1827] = -11'b00011010110; // -214
storage[1828] =  11'b00010010100; // 148
storage[1829] =  11'b00000110101; // 53
storage[1830] = -11'b00001011001; // -89
storage[1831] = -11'b00000110110; // -54
storage[1832] = -11'b00001001010; // -74
storage[1833] = -11'b00001001110; // -78
storage[1834] =  11'b00000110101; // 53
storage[1835] = -11'b00000101100; // -44
storage[1836] = -11'b00001100101; // -101
storage[1837] = -11'b00001011111; // -95
storage[1838] = -11'b00010000011; // -131
storage[1839] =  11'b00001000010; // 66
storage[1840] = -11'b00001110100; // -116
storage[1841] = -11'b00001110011; // -115
storage[1842] =  11'b00000010110; // 22
storage[1843] =  11'b00000110110; // 54
storage[1844] = -11'b00000000111; // -7
storage[1845] =  11'b00000101010; // 42
storage[1846] =  11'b00011001101; // 205
storage[1847] = -11'b00000111100; // -60
storage[1848] =  11'b00000001011; // 11
storage[1849] =  11'b00001101001; // 105
storage[1850] = -11'b00000011110; // -30
storage[1851] =  11'b00001100001; // 97
storage[1852] =  11'b00010000001; // 129
storage[1853] =  11'b00011011000; // 216
storage[1854] =  11'b00011010110; // 214
storage[1855] =  11'b00011000001; // 193
storage[1856] =  11'b00000011001; // 25
storage[1857] = -11'b00000011110; // -30
storage[1858] =  11'b00001111100; // 124
storage[1859] = -11'b00000110111; // -55
storage[1860] =  11'b00000001001; // 9
storage[1861] =  11'b00000101101; // 45
storage[1862] =  11'b00010000010; // 130
storage[1863] =  11'b00011000100; // 196
storage[1864] = -11'b00000011011; // -27
storage[1865] = -11'b00001111111; // -127
storage[1866] =  11'b00000000001; // 1
storage[1867] = -11'b00001011101; // -93
storage[1868] = -11'b00001100011; // -99
storage[1869] = -11'b00000010011; // -19
storage[1870] = -11'b00000011111; // -31
storage[1871] = -11'b00000011010; // -26
storage[1872] =  11'b00001111100; // 124
storage[1873] = -11'b00001101000; // -104
storage[1874] = -11'b00000000011; // -3
storage[1875] =  11'b00000101011; // 43
storage[1876] = -11'b00001101100; // -108
storage[1877] = -11'b00000110110; // -54
storage[1878] =  11'b00000010110; // 22
storage[1879] =  11'b00000001110; // 14
storage[1880] = -11'b00010010000; // -144
storage[1881] =  11'b00001011101; // 93
storage[1882] =  11'b00010011010; // 154
storage[1883] =  11'b00000110100; // 52
storage[1884] =  11'b00010001111; // 143
storage[1885] =  11'b00010011101; // 157
storage[1886] =  11'b00000110110; // 54
storage[1887] =  11'b00010000101; // 133
storage[1888] =  11'b00000011001; // 25
storage[1889] = -11'b00000001101; // -13
storage[1890] = -11'b00000001001; // -9
storage[1891] =  11'b00001001001; // 73
storage[1892] = -11'b00000110010; // -50
storage[1893] =  11'b00001111101; // 125
storage[1894] =  11'b00000101111; // 47
storage[1895] =  11'b00010000011; // 131
storage[1896] =  11'b00001000111; // 71
storage[1897] =  11'b00000101111; // 47
storage[1898] = -11'b00010001011; // -139
storage[1899] =  11'b00000001111; // 15
storage[1900] = -11'b00000001100; // -12
storage[1901] = -11'b00000010111; // -23
storage[1902] =  11'b00011001100; // 204
storage[1903] =  11'b00001010101; // 85
storage[1904] =  11'b00010111011; // 187
storage[1905] =  11'b00010010010; // 146
storage[1906] =  11'b00000101000; // 40
storage[1907] =  11'b00001011001; // 89
storage[1908] = -11'b00001001110; // -78
storage[1909] = -11'b00001001111; // -79
storage[1910] = -11'b00010000010; // -130
storage[1911] = -11'b00000000010; // -2
storage[1912] =  11'b00001000101; // 69
storage[1913] = -11'b00001101000; // -104
storage[1914] =  11'b00000110110; // 54
storage[1915] =  11'b00001011001; // 89
storage[1916] = -11'b00001010101; // -85
storage[1917] =  11'b00000011011; // 27
storage[1918] = -11'b00100011010; // -282
storage[1919] = -11'b00100100000; // -288
storage[1920] = -11'b00010111110; // -190
storage[1921] = -11'b00011000011; // -195
storage[1922] = -11'b00010001001; // -137
storage[1923] = -11'b00000000010; // -2
storage[1924] =  11'b00011000010; // 194
storage[1925] =  11'b00001111101; // 125
storage[1926] =  11'b00001001001; // 73
storage[1927] = -11'b00010011000; // -152
storage[1928] = -11'b00011010000; // -208
storage[1929] =  11'b00000111000; // 56
storage[1930] = -11'b00001010001; // -81
storage[1931] = -11'b00000010010; // -18
storage[1932] =  11'b00011000000; // 192
storage[1933] =  11'b00010110110; // 182
storage[1934] =  11'b00001001111; // 79
storage[1935] =  11'b00001010100; // 84
storage[1936] = -11'b00000000110; // -6
storage[1937] =  11'b00001000111; // 71
storage[1938] = -11'b00000010011; // -19
storage[1939] =  11'b00001100111; // 103
storage[1940] =  11'b00000111110; // 62
storage[1941] =  11'b00001001111; // 79
storage[1942] =  11'b00000110101; // 53
storage[1943] =  11'b00000001000; // 8
storage[1944] =  11'b00001010011; // 83
storage[1945] =  11'b00000010010; // 18
storage[1946] =  11'b00001011110; // 94
storage[1947] =  11'b00001101110; // 110
storage[1948] =  11'b00001001011; // 75
storage[1949] =  11'b00000100111; // 39
storage[1950] =  11'b00000001100; // 12
storage[1951] =  11'b00010010011; // 147
storage[1952] =  11'b00000010001; // 17
storage[1953] = -11'b00000100011; // -35
storage[1954] = -11'b00000001011; // -11
storage[1955] = -11'b00000110110; // -54
storage[1956] =  11'b00010001100; // 140
storage[1957] = -11'b00011011111; // -223
storage[1958] = -11'b00011100011; // -227
storage[1959] = -11'b00001001101; // -77
storage[1960] =  11'b00000001001; // 9
storage[1961] = -11'b00001011000; // -88
storage[1962] =  11'b00000001010; // 10
storage[1963] = -11'b00101010101; // -341
storage[1964] = -11'b00011100010; // -226
storage[1965] =  11'b00001110101; // 117
storage[1966] = -11'b00101100001; // -353
storage[1967] = -11'b00001100101; // -101
storage[1968] =  11'b00010000001; // 129
storage[1969] =  11'b00000000101; // 5
storage[1970] = -11'b00001000111; // -71
storage[1971] =  11'b00001001111; // 79
storage[1972] =  11'b00010110011; // 179
storage[1973] =  11'b00001110101; // 117
storage[1974] =  11'b00100001100; // 268
storage[1975] = -11'b00010001100; // -140
storage[1976] =  11'b00001000010; // 66
storage[1977] =  11'b00001110011; // 115
storage[1978] = -11'b00001111110; // -126
storage[1979] =  11'b00000100010; // 34
storage[1980] =  11'b00011001101; // 205
storage[1981] = -11'b00000001010; // -10
storage[1982] = -11'b00001001001; // -73
storage[1983] = -11'b00000001011; // -11
storage[1984] =  11'b00010000101; // 133
storage[1985] = -11'b00001000000; // -64
storage[1986] = -11'b00000011110; // -30
storage[1987] =  11'b00000101111; // 47
storage[1988] = -11'b00000010000; // -16
storage[1989] = -11'b00000111101; // -61
storage[1990] = -11'b00000110110; // -54
storage[1991] = -11'b00001000001; // -65
storage[1992] = -11'b00001010011; // -83
storage[1993] = -11'b00001010101; // -85
storage[1994] = -11'b00001101001; // -105
storage[1995] = -11'b00001001011; // -75
storage[1996] =  11'b00001110111; // 119
storage[1997] =  11'b00010101101; // 173
storage[1998] =  11'b00000110101; // 53
storage[1999] = -11'b00001110101; // -117
storage[2000] = -11'b00001010000; // -80
storage[2001] =  11'b00001110011; // 115
storage[2002] = -11'b00000011000; // -24
storage[2003] = -11'b00000010101; // -21
storage[2004] =  11'b00000101111; // 47
storage[2005] = -11'b00001010101; // -85
storage[2006] =  11'b00000110000; // 48
storage[2007] =  11'b00000111110; // 62
storage[2008] =  11'b00000011011; // 27
storage[2009] = -11'b00000001101; // -13
storage[2010] = -11'b00001110111; // -119
storage[2011] =  11'b00000100001; // 33
storage[2012] =  11'b00000100101; // 37
storage[2013] =  11'b00001100010; // 98
storage[2014] =  11'b00001110100; // 116
storage[2015] =  11'b00001110111; // 119
storage[2016] =  11'b00000000110; // 6
storage[2017] =  11'b00000001001; // 9
storage[2018] = -11'b00000101000; // -40
storage[2019] =  11'b00001111010; // 122
storage[2020] = -11'b00001000010; // -66
storage[2021] = -11'b00000100001; // -33
storage[2022] =  11'b00000110110; // 54
storage[2023] = -11'b00001011101; // -93
storage[2024] = -11'b00000101111; // -47
storage[2025] =  11'b00001011001; // 89
storage[2026] = -11'b00001101010; // -106
storage[2027] =  11'b00000010011; // 19
storage[2028] = -11'b00011011100; // -220
storage[2029] =  11'b00001101001; // 105
storage[2030] =  11'b00001111100; // 124
storage[2031] =  11'b00000111111; // 63
storage[2032] =  11'b00010011010; // 154
storage[2033] = -11'b00000100001; // -33
storage[2034] = -11'b00001100000; // -96
storage[2035] = -11'b00001000110; // -70
storage[2036] = -11'b00011101101; // -237
storage[2037] = -11'b00010011010; // -154
storage[2038] =  11'b00001101101; // 109
storage[2039] = -11'b00000001101; // -13
storage[2040] =  11'b00000111100; // 60
storage[2041] =  11'b00011011100; // 220
storage[2042] = -11'b00000010101; // -21
storage[2043] =  11'b00001011010; // 90
storage[2044] = -11'b00001000000; // -64
storage[2045] =  11'b00011111000; // 248
storage[2046] =  11'b00011001011; // 203
storage[2047] = -11'b00000011000; // -24
storage[2048] =  11'b00000011010; // 26
storage[2049] =  11'b00000000111; // 7
storage[2050] = -11'b00010010000; // -144
storage[2051] = -11'b00000010101; // -21
storage[2052] =  11'b00001100000; // 96
storage[2053] = -11'b00000011100; // -28
storage[2054] =  11'b00000001000; // 8
storage[2055] = -11'b00001111110; // -126
storage[2056] =  11'b00000001110; // 14
storage[2057] =  11'b00000010000; // 16
storage[2058] = -11'b00010100011; // -163
storage[2059] =  11'b00001000100; // 68
storage[2060] =  11'b00000110001; // 49
storage[2061] = -11'b00001110011; // -115
storage[2062] = -11'b00000111110; // -62
storage[2063] = -11'b00010011001; // -153
storage[2064] =  11'b00001000010; // 66
storage[2065] =  11'b00000111000; // 56
storage[2066] = -11'b00000000001; // -1
storage[2067] =  11'b00000101011; // 43
storage[2068] =  11'b00000010001; // 17
storage[2069] =  11'b00001001100; // 76
storage[2070] =  11'b00001101001; // 105
storage[2071] = -11'b00000000111; // -7
storage[2072] =  11'b00010010001; // 145
storage[2073] =  11'b00010101101; // 173
storage[2074] =  11'b00000100100; // 36
storage[2075] =  11'b00000101101; // 45
storage[2076] =  11'b00001001100; // 76
storage[2077] = -11'b00000010000; // -16
storage[2078] =  11'b00000101011; // 43
storage[2079] =  11'b00000001111; // 15
storage[2080] = -11'b00010000011; // -131
storage[2081] = -11'b00001101110; // -110
storage[2082] = -11'b00001110001; // -113
storage[2083] =  11'b00000011011; // 27
storage[2084] = -11'b00001001101; // -77
storage[2085] = -11'b00000010100; // -20
storage[2086] =  11'b00000100101; // 37
storage[2087] =  11'b00000001000; // 8
storage[2088] = -11'b00001001111; // -79
storage[2089] = -11'b00000100000; // -32
storage[2090] =  11'b00011001001; // 201
storage[2091] = -11'b00000010111; // -23
storage[2092] =  11'b00000010111; // 23
storage[2093] =  11'b00000111010; // 58
storage[2094] = -11'b00001110000; // -112
storage[2095] =  11'b00000101000; // 40
storage[2096] = -11'b00000110001; // -49
storage[2097] = -11'b00001100000; // -96
storage[2098] =  11'b00000001110; // 14
storage[2099] = -11'b00001001110; // -78
storage[2100] = -11'b00000100000; // -32
storage[2101] =  11'b00010011011; // 155
storage[2102] = -11'b00001101100; // -108
storage[2103] = -11'b00000101110; // -46
storage[2104] =  11'b00011001001; // 201
storage[2105] =  11'b00001011101; // 93
storage[2106] =  11'b00010100100; // 164
storage[2107] = -11'b00001110010; // -114
storage[2108] =  11'b00001010010; // 82
storage[2109] =  11'b00010011011; // 155
storage[2110] =  11'b00010001011; // 139
storage[2111] =  11'b00000101011; // 43
storage[2112] =  11'b00000011111; // 31
storage[2113] =  11'b00100000010; // 258
storage[2114] =  11'b00010100011; // 163
storage[2115] =  11'b00001010010; // 82
storage[2116] = -11'b00001111011; // -123
storage[2117] = -11'b00011011100; // -220
storage[2118] = -11'b00010000111; // -135
storage[2119] = -11'b00011100011; // -227
storage[2120] = -11'b00010100001; // -161
storage[2121] = -11'b00001001101; // -77
storage[2122] = -11'b00010011111; // -159
storage[2123] = -11'b00000101010; // -42
storage[2124] = -11'b00001011110; // -94
storage[2125] =  11'b00010110100; // 180
storage[2126] =  11'b00010000001; // 129
storage[2127] =  11'b00011011110; // 222
storage[2128] =  11'b00000110000; // 48
storage[2129] =  11'b00000000010; // 2
storage[2130] =  11'b00010000110; // 134
storage[2131] = -11'b00000001001; // -9
storage[2132] =  11'b00010010110; // 150
storage[2133] =  11'b00001111100; // 124
storage[2134] =  11'b00000010001; // 17
storage[2135] = -11'b00001011111; // -95
storage[2136] = -11'b00011011000; // -216
storage[2137] = -11'b00001000100; // -68
storage[2138] = -11'b00001101001; // -105
storage[2139] = -11'b00001001111; // -79
storage[2140] = -11'b00000111001; // -57
storage[2141] = -11'b00010010100; // -148
storage[2142] =  11'b00001010100; // 84
storage[2143] =  11'b00001010110; // 86
storage[2144] = -11'b00000100111; // -39
storage[2145] = -11'b00011010011; // -211
storage[2146] =  11'b00001000101; // 69
storage[2147] = -11'b00001111111; // -127
storage[2148] = -11'b00001001101; // -77
storage[2149] = -11'b00000111111; // -63
storage[2150] =  11'b00000110011; // 51
storage[2151] =  11'b00000101111; // 47
storage[2152] =  11'b00000011111; // 31
storage[2153] = -11'b00000100010; // -34
storage[2154] =  11'b00010011010; // 154
storage[2155] =  11'b00010000000; // 128
storage[2156] =  11'b00001000000; // 64
storage[2157] =  11'b00000011100; // 28
storage[2158] =  11'b00000110111; // 55
storage[2159] =  11'b00000010110; // 22
storage[2160] = -11'b00000110010; // -50
storage[2161] =  11'b00000100101; // 37
storage[2162] = -11'b00001011010; // -90
storage[2163] =  11'b00000111011; // 59
storage[2164] = -11'b00010001101; // -141
storage[2165] =  11'b00000000001; // 1
storage[2166] =  11'b00001101111; // 111
storage[2167] = -11'b00001011010; // -90
storage[2168] =  11'b00000010010; // 18
storage[2169] = -11'b00000101110; // -46
storage[2170] = -11'b00000001001; // -9
storage[2171] = -11'b00100101000; // -296
storage[2172] = -11'b00100111110; // -318
storage[2173] = -11'b00000101011; // -43
storage[2174] = -11'b00011000011; // -195
storage[2175] = -11'b00000111010; // -58
storage[2176] = -11'b00000010011; // -19
storage[2177] = -11'b00000111110; // -62
storage[2178] = -11'b00000000001; // -1
storage[2179] =  11'b00010101000; // 168
storage[2180] = -11'b00001000001; // -65
storage[2181] = -11'b00000001010; // -10
storage[2182] =  11'b00000110000; // 48
storage[2183] =  11'b00001111101; // 125
storage[2184] =  11'b00001010111; // 87
storage[2185] =  11'b00000111110; // 62
storage[2186] =  11'b00010111011; // 187
storage[2187] =  11'b00010011110; // 158
storage[2188] = -11'b00001011010; // -90
storage[2189] =  11'b00000110100; // 52
storage[2190] = -11'b00000010010; // -18
storage[2191] =  11'b00000111011; // 59
storage[2192] =  11'b00000010111; // 23
storage[2193] = -11'b00000001011; // -11
storage[2194] =  11'b00000111010; // 58
storage[2195] =  11'b00010101000; // 168
storage[2196] = -11'b00000011101; // -29
storage[2197] = -11'b00010000110; // -134
storage[2198] = -11'b00001011000; // -88
storage[2199] =  11'b00000001101; // 13
storage[2200] = -11'b00001000111; // -71
storage[2201] =  11'b00001001001; // 73
storage[2202] = -11'b00000101110; // -46
storage[2203] = -11'b00001001000; // -72
storage[2204] =  11'b00000110001; // 49
storage[2205] = -11'b00001000101; // -69
storage[2206] = -11'b00001000100; // -68
storage[2207] = -11'b00000010010; // -18
storage[2208] = -11'b00001111010; // -122
storage[2209] = -11'b00000000101; // -5
storage[2210] =  11'b00000100101; // 37
storage[2211] =  11'b00000110011; // 51
storage[2212] = -11'b00000001111; // -15
storage[2213] =  11'b00001111100; // 124
storage[2214] =  11'b00000100011; // 35
storage[2215] = -11'b00000011010; // -26
storage[2216] =  11'b00001000110; // 70
storage[2217] = -11'b00001111010; // -122
storage[2218] = -11'b00000101100; // -44
storage[2219] =  11'b00000101110; // 46
storage[2220] =  11'b00000101111; // 47
storage[2221] = -11'b00000000111; // -7
storage[2222] =  11'b00001000000; // 64
storage[2223] =  11'b00010000001; // 129
storage[2224] = -11'b00000111111; // -63
storage[2225] =  11'b00001111111; // 127
storage[2226] =  11'b00000001111; // 15
storage[2227] = -11'b00001100011; // -99
storage[2228] = -11'b00001101100; // -108
storage[2229] = -11'b00000010111; // -23
storage[2230] =  11'b00000110010; // 50
storage[2231] = -11'b00000110101; // -53
storage[2232] =  11'b00000110101; // 53
storage[2233] = -11'b00001101010; // -106
storage[2234] =  11'b00001111001; // 121
storage[2235] =  11'b00000110110; // 54
storage[2236] =  11'b00001000110; // 70
storage[2237] =  11'b00010000000; // 128
storage[2238] =  11'b00000111010; // 58
storage[2239] =  11'b00000101011; // 43
storage[2240] =  11'b00001000111; // 71
storage[2241] =  11'b00001010010; // 82
storage[2242] =  11'b00000011111; // 31
storage[2243] =  11'b00000010100; // 20
storage[2244] = -11'b00000110010; // -50
storage[2245] =  11'b00010010000; // 144
storage[2246] =  11'b00010110101; // 181
storage[2247] =  11'b00000011011; // 27
storage[2248] =  11'b00000100001; // 33
storage[2249] =  11'b00000000010; // 2
storage[2250] = -11'b00001100110; // -102
storage[2251] = -11'b00001011011; // -91
storage[2252] =  11'b00001101111; // 111
storage[2253] = -11'b00000110001; // -49
storage[2254] =  11'b00001110001; // 113
storage[2255] =  11'b00011010111; // 215
storage[2256] =  11'b00000011011; // 27
storage[2257] = -11'b00000001110; // -14
storage[2258] = -11'b00000100110; // -38
storage[2259] =  11'b00000011010; // 26
storage[2260] =  11'b00000000111; // 7
storage[2261] = -11'b00000000110; // -6
storage[2262] =  11'b00000110010; // 50
storage[2263] = -11'b00001011000; // -88
storage[2264] =  11'b00001001011; // 75
storage[2265] =  11'b00001101111; // 111
storage[2266] =  11'b00000110011; // 51
storage[2267] =  11'b00000010011; // 19
storage[2268] =  11'b00001011010; // 90
storage[2269] = -11'b00001001100; // -76
storage[2270] =  11'b00000100111; // 39
storage[2271] =  11'b00000101011; // 43
storage[2272] =  11'b00000100000; // 32
storage[2273] = -11'b00000100001; // -33
storage[2274] = -11'b00000010001; // -17
storage[2275] =  11'b00001100001; // 97
storage[2276] = -11'b00000100000; // -32
storage[2277] = -11'b00000001101; // -13
storage[2278] =  11'b00001100011; // 99
storage[2279] =  11'b00001100111; // 103
storage[2280] = -11'b00000100111; // -39
storage[2281] =  11'b00010011111; // 159
storage[2282] =  11'b00001100011; // 99
storage[2283] = -11'b00001101001; // -105
storage[2284] =  11'b00010111100; // 188
storage[2285] =  11'b00010000000; // 128
storage[2286] = -11'b00010010010; // -146
storage[2287] =  11'b00010011110; // 158
storage[2288] =  11'b00010111100; // 188
storage[2289] =  11'b00000101100; // 44
storage[2290] =  11'b00000101000; // 40
storage[2291] = -11'b00000001110; // -14
storage[2292] = -11'b00000101001; // -41
storage[2293] =  11'b00000010101; // 21
storage[2294] =  11'b00001001111; // 79
storage[2295] =  11'b00000100111; // 39
storage[2296] = -11'b00000100010; // -34
storage[2297] =  11'b00000100110; // 38
storage[2298] = -11'b00000111001; // -57
storage[2299] = -11'b00010001010; // -138
storage[2300] = -11'b00000110100; // -52
storage[2301] =  11'b00001011111; // 95
storage[2302] =  11'b00001000011; // 67
storage[2303] = -11'b00001111011; // -123
storage[2304] =  11'b00000100010; // 34
storage[2305] =  11'b00001000001; // 65
storage[2306] =  11'b00001011110; // 94
storage[2307] =  11'b00000110011; // 51
storage[2308] = -11'b00000101001; // -41
storage[2309] =  11'b00000001010; // 10
storage[2310] = -11'b00000010101; // -21
storage[2311] = -11'b00000101101; // -45
storage[2312] =  11'b00000011001; // 25
storage[2313] =  11'b00000000111; // 7
storage[2314] =  11'b00010001100; // 140
storage[2315] = -11'b00000010011; // -19
storage[2316] = -11'b00000111010; // -58
storage[2317] =  11'b00100000110; // 262
storage[2318] =  11'b00001110001; // 113
storage[2319] = -11'b00011010011; // -211
storage[2320] =  11'b00001011100; // 92
storage[2321] = -11'b00000100101; // -37
storage[2322] = -11'b00010011011; // -155
storage[2323] = -11'b00000110001; // -49
storage[2324] = -11'b00000011001; // -25
storage[2325] = -11'b00101010110; // -342
storage[2326] =  11'b00010011001; // 153
storage[2327] = -11'b00010111100; // -188
storage[2328] = -11'b00101011111; // -351
storage[2329] =  11'b00000101110; // 46
storage[2330] = -11'b00010110101; // -181
storage[2331] = -11'b00000010011; // -19
storage[2332] =  11'b00001011011; // 91
storage[2333] = -11'b00010101000; // -168
storage[2334] = -11'b00001110000; // -112
storage[2335] =  11'b00010010110; // 150
storage[2336] = -11'b00000111001; // -57
storage[2337] = -11'b00000001110; // -14
storage[2338] =  11'b00010111011; // 187
storage[2339] = -11'b00010010100; // -148
storage[2340] = -11'b00001100100; // -100
storage[2341] =  11'b00000011010; // 26
storage[2342] =  11'b00001100101; // 101
storage[2343] =  11'b00000011110; // 30
storage[2344] =  11'b00000110000; // 48
storage[2345] =  11'b00001110010; // 114
storage[2346] =  11'b00001011001; // 89
storage[2347] =  11'b00000011110; // 30
storage[2348] =  11'b00000000011; // 3
storage[2349] =  11'b00000110010; // 50
storage[2350] =  11'b00001111111; // 127
storage[2351] =  11'b00000110001; // 49
storage[2352] = -11'b00001100110; // -102
storage[2353] = -11'b00001000011; // -67
storage[2354] =  11'b00001011111; // 95
storage[2355] = -11'b00010100100; // -164
storage[2356] =  11'b00001001000; // 72
storage[2357] =  11'b00001111111; // 127
storage[2358] =  11'b00001011111; // 95
storage[2359] =  11'b00010001000; // 136
storage[2360] =  11'b00010110011; // 179
storage[2361] = -11'b00100110000; // -304
storage[2362] =  11'b00001001000; // 72
storage[2363] = -11'b00000100011; // -35
storage[2364] = -11'b00011111011; // -251
storage[2365] =  11'b00000101010; // 42
storage[2366] =  11'b00001000011; // 67
storage[2367] =  11'b00000011001; // 25
storage[2368] =  11'b00000011101; // 29
storage[2369] =  11'b00001001010; // 74
storage[2370] =  11'b00000010000; // 16
storage[2371] =  11'b00001100100; // 100
storage[2372] = -11'b00000110101; // -53
storage[2373] =  11'b00010010111; // 151
storage[2374] =  11'b00000000111; // 7
storage[2375] =  11'b00000100010; // 34
storage[2376] = -11'b00001011011; // -91
storage[2377] = -11'b00000000101; // -5
storage[2378] = -11'b00000010000; // -16
storage[2379] = -11'b00011101110; // -238
storage[2380] =  11'b00001100110; // 102
storage[2381] = -11'b00000000110; // -6
storage[2382] = -11'b00100011000; // -280
storage[2383] =  11'b00001001100; // 76
storage[2384] =  11'b00001111000; // 120
storage[2385] = -11'b00010101010; // -170
storage[2386] = -11'b00001000110; // -70
storage[2387] = -11'b00000011101; // -29
storage[2388] = -11'b00000110011; // -51
storage[2389] =  11'b00000000110; // 6
storage[2390] =  11'b00000000001; // 1
storage[2391] = -11'b00101110111; // -375
storage[2392] =  11'b00000000111; // 7
storage[2393] =  11'b00000001011; // 11
storage[2394] = -11'b00001000111; // -71
storage[2395] = -11'b00000100111; // -39
storage[2396] = -11'b00000011110; // -30
storage[2397] = -11'b00111010000; // -464
storage[2398] =  11'b00000101000; // 40
storage[2399] = -11'b00001111111; // -127
storage[2400] = -11'b00100101100; // -300
storage[2401] =  11'b00000001101; // 13
storage[2402] = -11'b00000001111; // -15
storage[2403] = -11'b00001100110; // -102
storage[2404] =  11'b00001000010; // 66
storage[2405] =  11'b00000111010; // 58
storage[2406] =  11'b00001011000; // 88
storage[2407] =  11'b00000110011; // 51
storage[2408] =  11'b00001001001; // 73
storage[2409] =  11'b00011000111; // 199
storage[2410] = -11'b00000101111; // -47
storage[2411] =  11'b00010010011; // 147
storage[2412] = -11'b00000100101; // -37
storage[2413] = -11'b00000110010; // -50
storage[2414] = -11'b00000011001; // -25
storage[2415] = -11'b00001001100; // -76
storage[2416] =  11'b00001000110; // 70
storage[2417] = -11'b00000011000; // -24
storage[2418] = -11'b00010001100; // -140
storage[2419] =  11'b00000010101; // 21
storage[2420] =  11'b00000100111; // 39
storage[2421] = -11'b00000001100; // -12
storage[2422] = -11'b00010001001; // -137
storage[2423] = -11'b00000010000; // -16
storage[2424] = -11'b00000101010; // -42
storage[2425] = -11'b00000111100; // -60
storage[2426] =  11'b00010001010; // 138
storage[2427] =  11'b00011000110; // 198
storage[2428] =  11'b00001011101; // 93
storage[2429] = -11'b00000011100; // -28
storage[2430] = -11'b00010001101; // -141
storage[2431] = -11'b00000010010; // -18
storage[2432] = -11'b00001111010; // -122
storage[2433] = -11'b00101100010; // -354
storage[2434] =  11'b00001010111; // 87
storage[2435] =  11'b00011010111; // 215
storage[2436] =  11'b00010111010; // 186
storage[2437] = -11'b00000000010; // -2
storage[2438] = -11'b00001000110; // -70
storage[2439] = -11'b00000011100; // -28
storage[2440] = -11'b00000000110; // -6
storage[2441] = -11'b00001100010; // -98
storage[2442] = -11'b00000110111; // -55
storage[2443] = -11'b00001110011; // -115
storage[2444] = -11'b00001000110; // -70
storage[2445] = -11'b00000010001; // -17
storage[2446] =  11'b00000011001; // 25
storage[2447] =  11'b00001101011; // 107
storage[2448] = -11'b00010001000; // -136
storage[2449] =  11'b00000000111; // 7
storage[2450] = -11'b00001000111; // -71
storage[2451] = -11'b00010001001; // -137
storage[2452] =  11'b00000100101; // 37
storage[2453] =  11'b00001011011; // 91
storage[2454] =  11'b00000011011; // 27
storage[2455] = -11'b00001011001; // -89
storage[2456] =  11'b00000101000; // 40
storage[2457] = -11'b00000111000; // -56
storage[2458] = -11'b00000110101; // -53
storage[2459] =  11'b00000111011; // 59
storage[2460] = -11'b00001011001; // -89
storage[2461] =  11'b00011010000; // 208
storage[2462] = -11'b00000001011; // -11
storage[2463] = -11'b00000110101; // -53
storage[2464] = -11'b00000010010; // -18
storage[2465] = -11'b00001000001; // -65
storage[2466] =  11'b00000110110; // 54
storage[2467] = -11'b00000010110; // -22
storage[2468] =  11'b00011000101; // 197
storage[2469] = -11'b00010101000; // -168
storage[2470] = -11'b00000000101; // -5
storage[2471] =  11'b00010000011; // 131
storage[2472] = -11'b00000001101; // -13
storage[2473] = -11'b00001100000; // -96
storage[2474] =  11'b00000100110; // 38
storage[2475] =  11'b00010111011; // 187
storage[2476] =  11'b00000100101; // 37
storage[2477] =  11'b00001101001; // 105
storage[2478] =  11'b00001000100; // 68
storage[2479] = -11'b00000001110; // -14
storage[2480] =  11'b00000011101; // 29
storage[2481] =  11'b00000110001; // 49
storage[2482] = -11'b00000110001; // -49
storage[2483] = -11'b00010011000; // -152
storage[2484] = -11'b00011001011; // -203
storage[2485] =  11'b00010000000; // 128
storage[2486] =  11'b00000110110; // 54
storage[2487] =  11'b00000001100; // 12
storage[2488] =  11'b00001010101; // 85
storage[2489] =  11'b00000010111; // 23
storage[2490] =  11'b00000000000; // 0
storage[2491] = -11'b00000011011; // -27
storage[2492] = -11'b00010011000; // -152
storage[2493] =  11'b00001000100; // 68
storage[2494] = -11'b00000110111; // -55
storage[2495] = -11'b00000011001; // -25
storage[2496] = -11'b00000101011; // -43
storage[2497] = -11'b00000011100; // -28
storage[2498] =  11'b00000100101; // 37
storage[2499] =  11'b00001010001; // 81
storage[2500] = -11'b00000100011; // -35
storage[2501] = -11'b00100000000; // -256
storage[2502] = -11'b00011000000; // -192
storage[2503] = -11'b00010010111; // -151
storage[2504] = -11'b00010011010; // -154
storage[2505] = -11'b00001011011; // -91
storage[2506] =  11'b00000011111; // 31
storage[2507] =  11'b00001100010; // 98
storage[2508] = -11'b00001111100; // -124
storage[2509] = -11'b00000001001; // -9
storage[2510] = -11'b00010011010; // -154
storage[2511] = -11'b00001101100; // -108
storage[2512] =  11'b00001010011; // 83
storage[2513] = -11'b00000001001; // -9
storage[2514] =  11'b00010001010; // 138
storage[2515] =  11'b00011011000; // 216
storage[2516] =  11'b00010010011; // 147
storage[2517] =  11'b00010111010; // 186
storage[2518] = -11'b00000000110; // -6
storage[2519] = -11'b00001001101; // -77
storage[2520] = -11'b00001001011; // -75
storage[2521] =  11'b00000001001; // 9
storage[2522] = -11'b00001110010; // -114
storage[2523] = -11'b00011001001; // -201
storage[2524] =  11'b00001101100; // 108
storage[2525] =  11'b00001100001; // 97
storage[2526] =  11'b00010001110; // 142
storage[2527] = -11'b00000000110; // -6
storage[2528] = -11'b00001010011; // -83
storage[2529] = -11'b00001101010; // -106
storage[2530] = -11'b00000101100; // -44
storage[2531] = -11'b00010000111; // -135
storage[2532] = -11'b00000011010; // -26
storage[2533] = -11'b00000111111; // -63
storage[2534] = -11'b00001000100; // -68
storage[2535] =  11'b00010110000; // 176
storage[2536] = -11'b00000101001; // -41
storage[2537] =  11'b00001000011; // 67
storage[2538] =  11'b00010011001; // 153
storage[2539] = -11'b00011010011; // -211
storage[2540] = -11'b00010010100; // -148
storage[2541] = -11'b00000101101; // -45
storage[2542] = -11'b00010110110; // -182
storage[2543] =  11'b00000011010; // 26
storage[2544] =  11'b00000001111; // 15
storage[2545] =  11'b00011010100; // 212
storage[2546] =  11'b00000101100; // 44
storage[2547] =  11'b00000100001; // 33
storage[2548] =  11'b00001001111; // 79
storage[2549] = -11'b00001001000; // -72
storage[2550] = -11'b00000010010; // -18
storage[2551] =  11'b00001000110; // 70
storage[2552] =  11'b00000011010; // 26
storage[2553] =  11'b00001011111; // 95
storage[2554] =  11'b00000101111; // 47
storage[2555] =  11'b00000000100; // 4
storage[2556] =  11'b00001001111; // 79
storage[2557] =  11'b00000111001; // 57
storage[2558] =  11'b00000101110; // 46
storage[2559] =  11'b00000101110; // 46
storage[2560] = -11'b00000001110; // -14
storage[2561] = -11'b00000001001; // -9
storage[2562] =  11'b00000110100; // 52
storage[2563] = -11'b00001101001; // -105
storage[2564] =  11'b00001010010; // 82
storage[2565] =  11'b00000100100; // 36
storage[2566] =  11'b00000101100; // 44
storage[2567] =  11'b00001110101; // 117
storage[2568] =  11'b00000001010; // 10
storage[2569] =  11'b00010100101; // 165
storage[2570] = -11'b00000110011; // -51
storage[2571] = -11'b00010011011; // -155
storage[2572] =  11'b00000000011; // 3
storage[2573] =  11'b00000010111; // 23
storage[2574] =  11'b00001011010; // 90
storage[2575] =  11'b00001011110; // 94
storage[2576] = -11'b00000000011; // -3
storage[2577] = -11'b00000011001; // -25
storage[2578] =  11'b00001111000; // 120
storage[2579] = -11'b00000011111; // -31
storage[2580] = -11'b00001010110; // -86
storage[2581] =  11'b00001011101; // 93
storage[2582] =  11'b00010010100; // 148
storage[2583] =  11'b00000100110; // 38
storage[2584] = -11'b00001100001; // -97
storage[2585] = -11'b00001010111; // -87
storage[2586] = -11'b00000101100; // -44
storage[2587] =  11'b00010000001; // 129
storage[2588] =  11'b00000010000; // 16
storage[2589] = -11'b00000101100; // -44
storage[2590] =  11'b00011010010; // 210
storage[2591] = -11'b00000100111; // -39
storage[2592] = -11'b00001101011; // -107
storage[2593] = -11'b00001011011; // -91
storage[2594] = -11'b00011110101; // -245
storage[2595] = -11'b00010101000; // -168
storage[2596] =  11'b00001001100; // 76
storage[2597] =  11'b00000001001; // 9
storage[2598] =  11'b00000010001; // 17
storage[2599] =  11'b00001001100; // 76
storage[2600] =  11'b00001101100; // 108
storage[2601] = -11'b00001100111; // -103
storage[2602] =  11'b00001111111; // 127
storage[2603] = -11'b00000000100; // -4
storage[2604] = -11'b00001010111; // -87
storage[2605] =  11'b00000011111; // 31
storage[2606] = -11'b00001001101; // -77
storage[2607] =  11'b00001111011; // 123
storage[2608] = -11'b00000110100; // -52
storage[2609] =  11'b00000011110; // 30
storage[2610] = -11'b00001011101; // -93
storage[2611] =  11'b00000000101; // 5
storage[2612] = -11'b00000111111; // -63
storage[2613] = -11'b00010010111; // -151
storage[2614] =  11'b00010000001; // 129
storage[2615] =  11'b00011111000; // 248
storage[2616] =  11'b00010000011; // 131
storage[2617] =  11'b00011110111; // 247
storage[2618] =  11'b00100000011; // 259
storage[2619] =  11'b00000000000; // 0
storage[2620] =  11'b00010010110; // 150
storage[2621] =  11'b00000000100; // 4
storage[2622] = -11'b00000011000; // -24
storage[2623] =  11'b00001011001; // 89
storage[2624] = -11'b00001001001; // -73
storage[2625] = -11'b00001111000; // -120
storage[2626] =  11'b00000001001; // 9
storage[2627] = -11'b00000101111; // -47
storage[2628] = -11'b00010011110; // -158
storage[2629] = -11'b00000111110; // -62
storage[2630] = -11'b00001100011; // -99
storage[2631] = -11'b00000110110; // -54
storage[2632] =  11'b00001001111; // 79
storage[2633] =  11'b00000011110; // 30
storage[2634] =  11'b00000100100; // 36
storage[2635] = -11'b00000000001; // -1
storage[2636] =  11'b00000001100; // 12
storage[2637] =  11'b00001011001; // 89
storage[2638] =  11'b00001111110; // 126
storage[2639] =  11'b00010010101; // 149
storage[2640] =  11'b00000100011; // 35
storage[2641] = -11'b00000101001; // -41
storage[2642] =  11'b00000010110; // 22
storage[2643] =  11'b00000111111; // 63
storage[2644] = -11'b00101100101; // -357
storage[2645] = -11'b00011000011; // -195
storage[2646] = -11'b00001111110; // -126
storage[2647] =  11'b00010000101; // 133
storage[2648] =  11'b00001010000; // 80
storage[2649] = -11'b00000011111; // -31
storage[2650] =  11'b00000110101; // 53
storage[2651] =  11'b00000001101; // 13
storage[2652] =  11'b00001011011; // 91
storage[2653] = -11'b00000000010; // -2
storage[2654] = -11'b00010000111; // -135
storage[2655] = -11'b00010001000; // -136
storage[2656] =  11'b00000000110; // 6
storage[2657] = -11'b00000100011; // -35
storage[2658] =  11'b00000111110; // 62
storage[2659] = -11'b00000011100; // -28
storage[2660] =  11'b00000001000; // 8
storage[2661] =  11'b00000101110; // 46
storage[2662] = -11'b00001110001; // -113
storage[2663] = -11'b00001011001; // -89
storage[2664] = -11'b00001010101; // -85
storage[2665] =  11'b00000110100; // 52
storage[2666] = -11'b00001101001; // -105
storage[2667] = -11'b00000110111; // -55
storage[2668] =  11'b00010101001; // 169
storage[2669] = -11'b00001100011; // -99
storage[2670] = -11'b00011011000; // -216
storage[2671] =  11'b00010101111; // 175
storage[2672] =  11'b00010011011; // 155
storage[2673] = -11'b00010000100; // -132
storage[2674] = -11'b00000101111; // -47
storage[2675] = -11'b00001100010; // -98
storage[2676] = -11'b00001110111; // -119
storage[2677] =  11'b00001110001; // 113
storage[2678] =  11'b00001110101; // 117
storage[2679] =  11'b00000001000; // 8
storage[2680] =  11'b00001110101; // 117
storage[2681] =  11'b00011011110; // 222
storage[2682] =  11'b00001110100; // 116
storage[2683] =  11'b00001010100; // 84
storage[2684] = -11'b00000011011; // -27
storage[2685] = -11'b00000101001; // -41
storage[2686] =  11'b00010000011; // 131
storage[2687] =  11'b00001110001; // 113
storage[2688] =  11'b00001110010; // 114
storage[2689] =  11'b00001111111; // 127
storage[2690] =  11'b00001010111; // 87
storage[2691] = -11'b00010000111; // -135
storage[2692] = -11'b00001010001; // -81
storage[2693] =  11'b00001101100; // 108
storage[2694] = -11'b00001110100; // -116
storage[2695] = -11'b00001101010; // -106
storage[2696] = -11'b00001010010; // -82
storage[2697] = -11'b00011110100; // -244
storage[2698] = -11'b00000110101; // -53
storage[2699] = -11'b00001000110; // -70
storage[2700] = -11'b00001101110; // -110
storage[2701] =  11'b00000011101; // 29
storage[2702] = -11'b00001100000; // -96
storage[2703] =  11'b00000110000; // 48
storage[2704] = -11'b00000001001; // -9
storage[2705] = -11'b00000101111; // -47
storage[2706] = -11'b00001001101; // -77
storage[2707] =  11'b00010111011; // 187
storage[2708] =  11'b00001100111; // 103
storage[2709] =  11'b00000101011; // 43
storage[2710] =  11'b00001010111; // 87
storage[2711] =  11'b00001000100; // 68
storage[2712] =  11'b00001110000; // 112
storage[2713] =  11'b00010100100; // 164
storage[2714] =  11'b00010111011; // 187
storage[2715] =  11'b00010001010; // 138
storage[2716] =  11'b00010000011; // 131
storage[2717] =  11'b00001001101; // 77
storage[2718] =  11'b00010011011; // 155
storage[2719] = -11'b00000100101; // -37
storage[2720] =  11'b00001101000; // 104
storage[2721] =  11'b00000101110; // 46
storage[2722] = -11'b00000000010; // -2
storage[2723] =  11'b00001001101; // 77
storage[2724] =  11'b00010011001; // 153
storage[2725] = -11'b00000010011; // -19
storage[2726] =  11'b00001000111; // 71
storage[2727] = -11'b00000110111; // -55
storage[2728] =  11'b00001000010; // 66
storage[2729] = -11'b00000100111; // -39
storage[2730] = -11'b00000100110; // -38
storage[2731] = -11'b00000001111; // -15
storage[2732] = -11'b00000010100; // -20
storage[2733] =  11'b00001101010; // 106
storage[2734] =  11'b00001101101; // 109
storage[2735] = -11'b00000010111; // -23
storage[2736] = -11'b00000101111; // -47
storage[2737] = -11'b00000110001; // -49
storage[2738] = -11'b00000111010; // -58
storage[2739] = -11'b00001111100; // -124
storage[2740] = -11'b00010110000; // -176
storage[2741] = -11'b00010011000; // -152
storage[2742] = -11'b00100001110; // -270
storage[2743] = -11'b00000101000; // -40
storage[2744] =  11'b00000110000; // 48
storage[2745] = -11'b00001001011; // -75
storage[2746] = -11'b00010001000; // -136
storage[2747] = -11'b00011110011; // -243
storage[2748] = -11'b00010010101; // -149
storage[2749] = -11'b00000101111; // -47
storage[2750] = -11'b00000011001; // -25
storage[2751] = -11'b00000101010; // -42
storage[2752] =  11'b00010110110; // 182
storage[2753] =  11'b00011100000; // 224
storage[2754] =  11'b00010110010; // 178
storage[2755] = -11'b00001101111; // -111
storage[2756] = -11'b00001101000; // -104
storage[2757] =  11'b00000000100; // 4
storage[2758] = -11'b00011011001; // -217
storage[2759] = -11'b00000100000; // -32
storage[2760] =  11'b00000101100; // 44
storage[2761] =  11'b00001111001; // 121
storage[2762] =  11'b00011100101; // 229
storage[2763] =  11'b00001100111; // 103
storage[2764] = -11'b00001100010; // -98
storage[2765] = -11'b00000101100; // -44
storage[2766] =  11'b00000001000; // 8
storage[2767] = -11'b00010110110; // -182
storage[2768] = -11'b00101101100; // -364
storage[2769] = -11'b00010100100; // -164
storage[2770] = -11'b00001111000; // -120
storage[2771] = -11'b00100010101; // -277
storage[2772] = -11'b00100101100; // -300
storage[2773] =  11'b00000111011; // 59
storage[2774] =  11'b00001001000; // 72
storage[2775] = -11'b00000001101; // -13
storage[2776] =  11'b00000010001; // 17
storage[2777] =  11'b00000110110; // 54
storage[2778] =  11'b00000011101; // 29
storage[2779] =  11'b00001010101; // 85
storage[2780] =  11'b00001110001; // 113
storage[2781] =  11'b00000010101; // 21
storage[2782] =  11'b00000111100; // 60
storage[2783] = -11'b00000110111; // -55
storage[2784] =  11'b00001101100; // 108
storage[2785] =  11'b00000001000; // 8
storage[2786] = -11'b00001011101; // -93
storage[2787] = -11'b00000000110; // -6
storage[2788] = -11'b00000001000; // -8
storage[2789] = -11'b00010100011; // -163
storage[2790] = -11'b00100000111; // -263
storage[2791] =  11'b00001011000; // 88
storage[2792] =  11'b00000110001; // 49
storage[2793] =  11'b00010010101; // 149
storage[2794] = -11'b00000100001; // -33
storage[2795] = -11'b00010010111; // -151
storage[2796] = -11'b00000111001; // -57
storage[2797] =  11'b00001010101; // 85
storage[2798] = -11'b00010110100; // -180
storage[2799] = -11'b00001101100; // -108
storage[2800] =  11'b00000100010; // 34
storage[2801] =  11'b00000101111; // 47
storage[2802] =  11'b00001101010; // 106
storage[2803] =  11'b00001001000; // 72
storage[2804] = -11'b00000101101; // -45
storage[2805] = -11'b00001100101; // -101
storage[2806] = -11'b00000101101; // -45
storage[2807] = -11'b00000101010; // -42
storage[2808] =  11'b00000100110; // 38
storage[2809] =  11'b00000100011; // 35
storage[2810] =  11'b00001100111; // 103
storage[2811] =  11'b00000000101; // 5
storage[2812] =  11'b00000010000; // 16
storage[2813] =  11'b00001010000; // 80
storage[2814] = -11'b00000110001; // -49
storage[2815] = -11'b00000000001; // -1
storage[2816] = -11'b00001001100; // -76
storage[2817] = -11'b00001011110; // -94
storage[2818] =  11'b00000111101; // 61
storage[2819] = -11'b00000111000; // -56
storage[2820] =  11'b00001000000; // 64
storage[2821] =  11'b00001010110; // 86
storage[2822] =  11'b00010011110; // 158
storage[2823] =  11'b00001001111; // 79
storage[2824] = -11'b00000100111; // -39
storage[2825] =  11'b00000000001; // 1
storage[2826] =  11'b00010110000; // 176
storage[2827] =  11'b00000110110; // 54
storage[2828] = -11'b00000001010; // -10
storage[2829] =  11'b00001110101; // 117
storage[2830] =  11'b00000000100; // 4
storage[2831] =  11'b00001010111; // 87
storage[2832] = -11'b00001010000; // -80
storage[2833] =  11'b00001010101; // 85
storage[2834] =  11'b00001000000; // 64
storage[2835] = -11'b00001111110; // -126
storage[2836] =  11'b00011100110; // 230
storage[2837] =  11'b00001111010; // 122
storage[2838] =  11'b00001011110; // 94
storage[2839] =  11'b00000011010; // 26
storage[2840] =  11'b00000000010; // 2
storage[2841] =  11'b00000100101; // 37
storage[2842] =  11'b00000100000; // 32
storage[2843] = -11'b00010000111; // -135
storage[2844] =  11'b00000001100; // 12
storage[2845] =  11'b00010100101; // 165
storage[2846] =  11'b00000011000; // 24
storage[2847] =  11'b00000110101; // 53
storage[2848] =  11'b00001010010; // 82
storage[2849] = -11'b00000110111; // -55
storage[2850] =  11'b00001010011; // 83
storage[2851] = -11'b00000001101; // -13
storage[2852] =  11'b00000101010; // 42
storage[2853] =  11'b00011101010; // 234
storage[2854] =  11'b00001001011; // 75
storage[2855] = -11'b00010001010; // -138
storage[2856] = -11'b00000111000; // -56
storage[2857] =  11'b00001001100; // 76
storage[2858] = -11'b00011011010; // -218
storage[2859] = -11'b00000011110; // -30
storage[2860] = -11'b00001101101; // -109
storage[2861] = -11'b00001010000; // -80
storage[2862] =  11'b00001100101; // 101
storage[2863] =  11'b00000111000; // 56
storage[2864] = -11'b00000101101; // -45
storage[2865] =  11'b00001110000; // 112
storage[2866] =  11'b00001011011; // 91
storage[2867] = -11'b00010001100; // -140
storage[2868] = -11'b00001000100; // -68
storage[2869] =  11'b00000000110; // 6
storage[2870] = -11'b00000000011; // -3
storage[2871] =  11'b00000000010; // 2
storage[2872] = -11'b00001000100; // -68
storage[2873] = -11'b00010000101; // -133
storage[2874] = -11'b00000111111; // -63
storage[2875] = -11'b00000111111; // -63
storage[2876] =  11'b00000011110; // 30
storage[2877] = -11'b00000100011; // -35
storage[2878] =  11'b00000111011; // 59
storage[2879] =  11'b00001000011; // 67
storage[2880] = -11'b00000001111; // -15
storage[2881] =  11'b00011001111; // 207
storage[2882] =  11'b00001110101; // 117
storage[2883] =  11'b00000001110; // 14
storage[2884] =  11'b00010000001; // 129
storage[2885] = -11'b00010010001; // -145
storage[2886] = -11'b00000110110; // -54
storage[2887] = -11'b00000101111; // -47
storage[2888] =  11'b00000101000; // 40
storage[2889] =  11'b00000101100; // 44
storage[2890] =  11'b00001111111; // 127
storage[2891] =  11'b00100101101; // 301
storage[2892] =  11'b00001111001; // 121
storage[2893] =  11'b00000010011; // 19
storage[2894] = -11'b00011011100; // -220
storage[2895] = -11'b00000011010; // -26
storage[2896] = -11'b00001011100; // -92
storage[2897] =  11'b00000001110; // 14
storage[2898] =  11'b00000011011; // 27
storage[2899] =  11'b00011000011; // 195
storage[2900] = -11'b00000001001; // -9
storage[2901] = -11'b00000000101; // -5
storage[2902] = -11'b00010001110; // -142
storage[2903] = -11'b00100110110; // -310
storage[2904] = -11'b00000100111; // -39
storage[2905] = -11'b00001111101; // -125
storage[2906] = -11'b00000111000; // -56
storage[2907] = -11'b00001111101; // -125
storage[2908] =  11'b00001001100; // 76
storage[2909] = -11'b00000110001; // -49
storage[2910] =  11'b00000001011; // 11
storage[2911] = -11'b00001001110; // -78
storage[2912] = -11'b00001000001; // -65
storage[2913] = -11'b00000100101; // -37
storage[2914] =  11'b00001011101; // 93
storage[2915] =  11'b00000100101; // 37
storage[2916] =  11'b00001010100; // 84
storage[2917] =  11'b00001000010; // 66
storage[2918] = -11'b00000001000; // -8
storage[2919] =  11'b00000000111; // 7
storage[2920] =  11'b00000001110; // 14
storage[2921] =  11'b00000110010; // 50
storage[2922] = -11'b00000011011; // -27
storage[2923] = -11'b00000011111; // -31
storage[2924] =  11'b00000100011; // 35
storage[2925] = -11'b00000001110; // -14
storage[2926] =  11'b00001101000; // 104
storage[2927] =  11'b00000000100; // 4
storage[2928] =  11'b00000101100; // 44
storage[2929] =  11'b00001011000; // 88
storage[2930] =  11'b00000000101; // 5
storage[2931] =  11'b00000100010; // 34
storage[2932] =  11'b00000110011; // 51
storage[2933] =  11'b00001011000; // 88
storage[2934] = -11'b00001100010; // -98
storage[2935] =  11'b00001010001; // 81
storage[2936] =  11'b00000000001; // 1
storage[2937] =  11'b00001111111; // 127
storage[2938] =  11'b00001011000; // 88
storage[2939] = -11'b00001011010; // -90
storage[2940] =  11'b00000101010; // 42
storage[2941] = -11'b00000001111; // -15
storage[2942] =  11'b00000010110; // 22
storage[2943] = -11'b00000100101; // -37
storage[2944] = -11'b00001000111; // -71
storage[2945] = -11'b00010000101; // -133
storage[2946] = -11'b00000101011; // -43
storage[2947] = -11'b00000011010; // -26
storage[2948] = -11'b00000100101; // -37
storage[2949] = -11'b00000010111; // -23
storage[2950] = -11'b00010010101; // -149
storage[2951] = -11'b00001100011; // -99
storage[2952] = -11'b00010010110; // -150
storage[2953] =  11'b00001001010; // 74
storage[2954] =  11'b00000010000; // 16
storage[2955] = -11'b00000101001; // -41
storage[2956] =  11'b00001010010; // 82
storage[2957] = -11'b00000110101; // -53
storage[2958] =  11'b00000110100; // 52
storage[2959] = -11'b00000101111; // -47
storage[2960] = -11'b00000111011; // -59
storage[2961] =  11'b00010001111; // 143
storage[2962] = -11'b00000001101; // -13
storage[2963] =  11'b00001111111; // 127
storage[2964] =  11'b00000010011; // 19
storage[2965] =  11'b00000010101; // 21
storage[2966] =  11'b00010001011; // 139
storage[2967] =  11'b00011011001; // 217
storage[2968] = -11'b00001011000; // -88
storage[2969] =  11'b00010011100; // 156
storage[2970] =  11'b00010001010; // 138
storage[2971] =  11'b00001101111; // 111
storage[2972] =  11'b00100000001; // 257
storage[2973] =  11'b00001011101; // 93
storage[2974] =  11'b00011011100; // 220
storage[2975] =  11'b00011100110; // 230
storage[2976] =  11'b00011111111; // 255
storage[2977] = -11'b00000101111; // -47
storage[2978] =  11'b00010111000; // 184
storage[2979] =  11'b00001010101; // 85
storage[2980] = -11'b00000111110; // -62
storage[2981] = -11'b00000100010; // -34
storage[2982] = -11'b00001110100; // -116
storage[2983] =  11'b00001000110; // 70
storage[2984] = -11'b00000010000; // -16
storage[2985] = -11'b00001100010; // -98
storage[2986] =  11'b00001100010; // 98
storage[2987] =  11'b00000101001; // 41
storage[2988] = -11'b00001010101; // -85
storage[2989] = -11'b00001000100; // -68
storage[2990] =  11'b00000010100; // 20
storage[2991] =  11'b00000101000; // 40
storage[2992] =  11'b00000001010; // 10
storage[2993] =  11'b00000111000; // 56
storage[2994] =  11'b00000001101; // 13
storage[2995] =  11'b00000101010; // 42
storage[2996] = -11'b00000100001; // -33
storage[2997] =  11'b00000111111; // 63
storage[2998] =  11'b00001010001; // 81
storage[2999] =  11'b00000101111; // 47
storage[3000] =  11'b00000000110; // 6
storage[3001] =  11'b00000100010; // 34
storage[3002] =  11'b00000001001; // 9
storage[3003] = -11'b00000000101; // -5
storage[3004] = -11'b00000011111; // -31
storage[3005] = -11'b00000011111; // -31
storage[3006] = -11'b00010111000; // -184
storage[3007] = -11'b00000100110; // -38
storage[3008] = -11'b00000000100; // -4
storage[3009] = -11'b00000000110; // -6
storage[3010] =  11'b00000001101; // 13
storage[3011] =  11'b00000011010; // 26
storage[3012] = -11'b00001010000; // -80
storage[3013] =  11'b00000011001; // 25
storage[3014] =  11'b00001000001; // 65
storage[3015] = -11'b00001110000; // -112
storage[3016] =  11'b00001010011; // 83
storage[3017] =  11'b00001010001; // 81
storage[3018] =  11'b00000011100; // 28
storage[3019] =  11'b00001001111; // 79
storage[3020] =  11'b00000100110; // 38
storage[3021] =  11'b00001001000; // 72
storage[3022] =  11'b00001000111; // 71
storage[3023] =  11'b00000111100; // 60
storage[3024] =  11'b00001000001; // 65
storage[3025] = -11'b00000000001; // -1
storage[3026] = -11'b00000001010; // -10
storage[3027] = -11'b00000011010; // -26
storage[3028] =  11'b00000101000; // 40
storage[3029] = -11'b00000011000; // -24
storage[3030] = -11'b00001110111; // -119
storage[3031] = -11'b00000010100; // -20
storage[3032] = -11'b00000110111; // -55
storage[3033] = -11'b00011001011; // -203
storage[3034] = -11'b00001000001; // -65
storage[3035] = -11'b00000111000; // -56
storage[3036] = -11'b00000111100; // -60
storage[3037] = -11'b00001000010; // -66
storage[3038] =  11'b00000001010; // 10
storage[3039] =  11'b00000111010; // 58
storage[3040] =  11'b00000110101; // 53
storage[3041] =  11'b00001001011; // 75
storage[3042] =  11'b00000111101; // 61
storage[3043] = -11'b00000100001; // -33
storage[3044] =  11'b00000001101; // 13
storage[3045] =  11'b00000001111; // 15
storage[3046] = -11'b00000111011; // -59
storage[3047] =  11'b00000100101; // 37
storage[3048] =  11'b00001000101; // 69
storage[3049] = -11'b00001011010; // -90
storage[3050] =  11'b00000101110; // 46
storage[3051] =  11'b00001000101; // 69
storage[3052] = -11'b00001100100; // -100
storage[3053] =  11'b00000010000; // 16
storage[3054] =  11'b00000000000; // 0
storage[3055] = -11'b00000001001; // -9
storage[3056] =  11'b00000001100; // 12
storage[3057] =  11'b00000100011; // 35
storage[3058] = -11'b00000000011; // -3
storage[3059] =  11'b00000000110; // 6
storage[3060] =  11'b00000011111; // 31
storage[3061] =  11'b00000010101; // 21
storage[3062] = -11'b00000000001; // -1
storage[3063] =  11'b00000010000; // 16
storage[3064] = -11'b00000011000; // -24
storage[3065] =  11'b00000010010; // 18
storage[3066] =  11'b00010011000; // 152
storage[3067] = -11'b00000110101; // -53
storage[3068] =  11'b00000011001; // 25
storage[3069] = -11'b00010010010; // -146
storage[3070] =  11'b00000100001; // 33
storage[3071] = -11'b00000000111; // -7
storage[3072] = -11'b00000100110; // -38
storage[3073] =  11'b00001011010; // 90
storage[3074] =  11'b00000011000; // 24
storage[3075] =  11'b00000001110; // 14
storage[3076] =  11'b00000110011; // 51
storage[3077] = -11'b00000000111; // -7
storage[3078] = -11'b00000100011; // -35
storage[3079] = -11'b00010001010; // -138
storage[3080] = -11'b00000101111; // -47
storage[3081] =  11'b00000100010; // 34
storage[3082] = -11'b00010001110; // -142
storage[3083] = -11'b00001010100; // -84
storage[3084] = -11'b00000100111; // -39
storage[3085] =  11'b00000011001; // 25
storage[3086] = -11'b00000110010; // -50
storage[3087] = -11'b00001001000; // -72
storage[3088] =  11'b00000001101; // 13
storage[3089] =  11'b00000110000; // 48
storage[3090] = -11'b00000101101; // -45
storage[3091] = -11'b00000111011; // -59
storage[3092] = -11'b00000110011; // -51
storage[3093] = -11'b00010000010; // -130
storage[3094] = -11'b00000111110; // -62
storage[3095] = -11'b00001011001; // -89
storage[3096] = -11'b00001010100; // -84
storage[3097] = -11'b00000010100; // -20
storage[3098] = -11'b00000000111; // -7
storage[3099] = -11'b00000000100; // -4
storage[3100] = -11'b00000011001; // -25
storage[3101] =  11'b00000110110; // 54
storage[3102] = -11'b00000001111; // -15
storage[3103] = -11'b00001000000; // -64
storage[3104] = -11'b00000011010; // -26
storage[3105] =  11'b00000010110; // 22
storage[3106] = -11'b00010001011; // -139
storage[3107] =  11'b00001001110; // 78
storage[3108] =  11'b00000110011; // 51
storage[3109] =  11'b00000100011; // 35
storage[3110] =  11'b00000101011; // 43
storage[3111] =  11'b00000110001; // 49
storage[3112] =  11'b00001011000; // 88
storage[3113] = -11'b00000000100; // -4
storage[3114] =  11'b00000010111; // 23
storage[3115] = -11'b00000101011; // -43
storage[3116] = -11'b00001110010; // -114
storage[3117] = -11'b00011001101; // -205
storage[3118] =  11'b00000111111; // 63
storage[3119] =  11'b00000110010; // 50
storage[3120] = -11'b00000011111; // -31
storage[3121] =  11'b00000000011; // 3
storage[3122] = -11'b00000011011; // -27
storage[3123] = -11'b00000001100; // -12
storage[3124] = -11'b00000011000; // -24
storage[3125] =  11'b00000111110; // 62
storage[3126] =  11'b00001010010; // 82
storage[3127] =  11'b00000101010; // 42
storage[3128] =  11'b00000111110; // 62
storage[3129] =  11'b00000110011; // 51
storage[3130] =  11'b00000001101; // 13
storage[3131] =  11'b00000101100; // 44
storage[3132] =  11'b00000010010; // 18
storage[3133] =  11'b00000010001; // 17
storage[3134] = -11'b00000111100; // -60
storage[3135] = -11'b00000101111; // -47
storage[3136] = -11'b00000011111; // -31
storage[3137] =  11'b00000010110; // 22
storage[3138] = -11'b00000010101; // -21
storage[3139] =  11'b00000001101; // 13
storage[3140] = -11'b00000011101; // -29
storage[3141] =  11'b00000001010; // 10
storage[3142] =  11'b00000101010; // 42
storage[3143] =  11'b00000010000; // 16
storage[3144] = -11'b00000101000; // -40
storage[3145] = -11'b00000101111; // -47
storage[3146] = -11'b00001110001; // -113
storage[3147] = -11'b00001001101; // -77
storage[3148] =  11'b00000000001; // 1
storage[3149] = -11'b00000101010; // -42
storage[3150] = -11'b00000011010; // -26
storage[3151] =  11'b00000100011; // 35
storage[3152] =  11'b00000010110; // 22
storage[3153] = -11'b00000011011; // -27
storage[3154] = -11'b00000000111; // -7
storage[3155] =  11'b00000111100; // 60
storage[3156] =  11'b00000111001; // 57
storage[3157] =  11'b00000010001; // 17
storage[3158] = -11'b00000010001; // -17
storage[3159] =  11'b00000001001; // 9
storage[3160] = -11'b00001101010; // -106
storage[3161] =  11'b00000010011; // 19
storage[3162] = -11'b00000000111; // -7
storage[3163] = -11'b00000100000; // -32
storage[3164] =  11'b00000010001; // 17
storage[3165] = -11'b00000110100; // -52
storage[3166] =  11'b00001100100; // 100
storage[3167] = -11'b00001010001; // -81
storage[3168] = -11'b00000000101; // -5
storage[3169] = -11'b00000010110; // -22
storage[3170] =  11'b00000110000; // 48
storage[3171] =  11'b00000100000; // 32
storage[3172] =  11'b00000100000; // 32
storage[3173] =  11'b00000110101; // 53
storage[3174] =  11'b00001100010; // 98
storage[3175] =  11'b00000100100; // 36
storage[3176] =  11'b00000110100; // 52
storage[3177] = -11'b00000000100; // -4
storage[3178] =  11'b00000111110; // 62
storage[3179] = -11'b00001110001; // -113
storage[3180] =  11'b00000001001; // 9
storage[3181] =  11'b00000001001; // 9
storage[3182] = -11'b00000010110; // -22
storage[3183] = -11'b00000001001; // -9
storage[3184] =  11'b00000110111; // 55
storage[3185] =  11'b00001010010; // 82
storage[3186] =  11'b00000001011; // 11
storage[3187] = -11'b00000001110; // -14
storage[3188] = -11'b00010101011; // -171
storage[3189] =  11'b00000111010; // 58
storage[3190] = -11'b00001100011; // -99
storage[3191] = -11'b00001010010; // -82
storage[3192] =  11'b00000111111; // 63
storage[3193] = -11'b00000001010; // -10
storage[3194] =  11'b00000110000; // 48
storage[3195] = -11'b00000001101; // -13
storage[3196] =  11'b00000000101; // 5
storage[3197] =  11'b00000000010; // 2
storage[3198] = -11'b00000101100; // -44
storage[3199] = -11'b00000011011; // -27
storage[3200] = -11'b00000110110; // -54
storage[3201] =  11'b00010110100; // 180
storage[3202] = -11'b00001010110; // -86
storage[3203] = -11'b00000100100; // -36
storage[3204] =  11'b00001101101; // 109
storage[3205] = -11'b00000110011; // -51
storage[3206] = -11'b00000110000; // -48
storage[3207] =  11'b00000100000; // 32
storage[3208] = -11'b00000001011; // -11
storage[3209] = -11'b00001001010; // -74
storage[3210] = -11'b00001100001; // -97
storage[3211] =  11'b00000010010; // 18
storage[3212] = -11'b00001101111; // -111
storage[3213] =  11'b00000101011; // 43
storage[3214] =  11'b00001010011; // 83
storage[3215] =  11'b00000110011; // 51
storage[3216] =  11'b00000010000; // 16
storage[3217] = -11'b00000000010; // -2
storage[3218] = -11'b00000010000; // -16
storage[3219] = -11'b00000110111; // -55
storage[3220] = -11'b00000100111; // -39
storage[3221] = -11'b00000010101; // -21
storage[3222] =  11'b00000000111; // 7
storage[3223] =  11'b00000100001; // 33
storage[3224] = -11'b00000100100; // -36
storage[3225] = -11'b00001001001; // -73
storage[3226] =  11'b00000000101; // 5
storage[3227] =  11'b00000100010; // 34
storage[3228] = -11'b00000111101; // -61
storage[3229] = -11'b00001001000; // -72
storage[3230] =  11'b00000011000; // 24
storage[3231] =  11'b00000101110; // 46
storage[3232] =  11'b00000010111; // 23
storage[3233] =  11'b00001001101; // 77
storage[3234] = -11'b00000100000; // -32
storage[3235] = -11'b00000001010; // -10
storage[3236] = -11'b00000011101; // -29
storage[3237] = -11'b00001010011; // -83
storage[3238] =  11'b00001100001; // 97
storage[3239] =  11'b00001000110; // 70
storage[3240] =  11'b00000110110; // 54
storage[3241] =  11'b00001010110; // 86
storage[3242] = -11'b00000100100; // -36
storage[3243] = -11'b00000100111; // -39
storage[3244] =  11'b00000010001; // 17
storage[3245] = -11'b00000010111; // -23
storage[3246] = -11'b00000110000; // -48
storage[3247] = -11'b00000101100; // -44
storage[3248] = -11'b00000101010; // -42
storage[3249] =  11'b00000110100; // 52
storage[3250] =  11'b00000010111; // 23
storage[3251] = -11'b00000101000; // -40
storage[3252] = -11'b00001011001; // -89
storage[3253] =  11'b00000011110; // 30
storage[3254] = -11'b00000000010; // -2
storage[3255] =  11'b00000011011; // 27
storage[3256] =  11'b00000010101; // 21
storage[3257] = -11'b00000010101; // -21
storage[3258] = -11'b00001001000; // -72
storage[3259] =  11'b00000000101; // 5
storage[3260] =  11'b00000110001; // 49
storage[3261] =  11'b00000001101; // 13
storage[3262] =  11'b00000101011; // 43
storage[3263] = -11'b00000011110; // -30
storage[3264] =  11'b00000011011; // 27
storage[3265] =  11'b00000011010; // 26
storage[3266] = -11'b00000010000; // -16
storage[3267] =  11'b00000101101; // 45
storage[3268] = -11'b00000001110; // -14
storage[3269] = -11'b00000001010; // -10
storage[3270] = -11'b00011000101; // -197
storage[3271] = -11'b00000010000; // -16
storage[3272] = -11'b00000111000; // -56
storage[3273] = -11'b00001111100; // -124
storage[3274] = -11'b00001100111; // -103
storage[3275] = -11'b00001001010; // -74
storage[3276] =  11'b00001000100; // 68
storage[3277] = -11'b00010001110; // -142
storage[3278] = -11'b00000010011; // -19
storage[3279] = -11'b00001100110; // -102
storage[3280] = -11'b00010111110; // -190
storage[3281] = -11'b00001110100; // -116
storage[3282] = -11'b00000011001; // -25
storage[3283] = -11'b00001101111; // -111
storage[3284] =  11'b00000000010; // 2
storage[3285] =  11'b00000011101; // 29
storage[3286] =  11'b00001010111; // 87
storage[3287] =  11'b00000010011; // 19
storage[3288] =  11'b00000001000; // 8
storage[3289] = -11'b00000100010; // -34
storage[3290] = -11'b00001001111; // -79
storage[3291] =  11'b00000001001; // 9
storage[3292] = -11'b00010011110; // -158
storage[3293] = -11'b00000101101; // -45
storage[3294] =  11'b00000011000; // 24
storage[3295] = -11'b00000101000; // -40
storage[3296] = -11'b00001010110; // -86
storage[3297] = -11'b00001100001; // -97
storage[3298] = -11'b00000011101; // -29
storage[3299] = -11'b00001010110; // -86
storage[3300] = -11'b00001100101; // -101
storage[3301] = -11'b00000111110; // -62
storage[3302] = -11'b00010011000; // -152
storage[3303] = -11'b00000010101; // -21
storage[3304] =  11'b00000100011; // 35
storage[3305] =  11'b00000100011; // 35
storage[3306] =  11'b00000100000; // 32
storage[3307] = -11'b00000001010; // -10
storage[3308] =  11'b00000011001; // 25
storage[3309] = -11'b00000000100; // -4
storage[3310] =  11'b00000101010; // 42
storage[3311] = -11'b00000011011; // -27
storage[3312] =  11'b00000100010; // 34
storage[3313] = -11'b00000001110; // -14
storage[3314] = -11'b00000100011; // -35
storage[3315] = -11'b00000100110; // -38
storage[3316] =  11'b00000111000; // 56
storage[3317] = -11'b00000101101; // -45
storage[3318] =  11'b00000001011; // 11
storage[3319] = -11'b00000100111; // -39
storage[3320] =  11'b00000010111; // 23
storage[3321] =  11'b00000000110; // 6
storage[3322] =  11'b00000000001; // 1
storage[3323] =  11'b00000111011; // 59
storage[3324] = -11'b00000110001; // -49
storage[3325] =  11'b00000110010; // 50
storage[3326] =  11'b00000100001; // 33
storage[3327] = -11'b00000110100; // -52
storage[3328] = -11'b00001010101; // -85
storage[3329] = -11'b00001011011; // -91
storage[3330] =  11'b00000011000; // 24
storage[3331] =  11'b00000001110; // 14
storage[3332] = -11'b00000010110; // -22
storage[3333] =  11'b00000000001; // 1
storage[3334] =  11'b00000100001; // 33
storage[3335] = -11'b00001001000; // -72
storage[3336] = -11'b00000010101; // -21
storage[3337] = -11'b00001100001; // -97
storage[3338] = -11'b00001011101; // -93
storage[3339] =  11'b00000101100; // 44
storage[3340] = -11'b00001110101; // -117
storage[3341] = -11'b00010100111; // -167
storage[3342] = -11'b00000010101; // -21
storage[3343] = -11'b00000100110; // -38
storage[3344] = -11'b00001101111; // -111
storage[3345] = -11'b00000111110; // -62
storage[3346] = -11'b00011101100; // -236
storage[3347] = -11'b00010001110; // -142
storage[3348] = -11'b00000011010; // -26
storage[3349] = -11'b00011110110; // -246
storage[3350] = -11'b00000110000; // -48
storage[3351] =  11'b00000001101; // 13
storage[3352] = -11'b00001110100; // -116
storage[3353] = -11'b00001001100; // -76
storage[3354] = -11'b00000010111; // -23
storage[3355] = -11'b00000110100; // -52
storage[3356] = -11'b00000000110; // -6
storage[3357] =  11'b00000110010; // 50
storage[3358] =  11'b00001010011; // 83
storage[3359] =  11'b00000000111; // 7
storage[3360] = -11'b00000101101; // -45
storage[3361] =  11'b00000110111; // 55
storage[3362] = -11'b00000110111; // -55
storage[3363] = -11'b00000011100; // -28
storage[3364] = -11'b00001100000; // -96
storage[3365] = -11'b00010000101; // -133
storage[3366] = -11'b00000101101; // -45
storage[3367] =  11'b00000101011; // 43
storage[3368] =  11'b00000001011; // 11
storage[3369] =  11'b00000100111; // 39
storage[3370] =  11'b00000101000; // 40
storage[3371] = -11'b00000010011; // -19
storage[3372] = -11'b00000001001; // -9
storage[3373] =  11'b00000111001; // 57
storage[3374] = -11'b00010110010; // -178
storage[3375] =  11'b00000000100; // 4
storage[3376] =  11'b00000011100; // 28
storage[3377] = -11'b00000000111; // -7
storage[3378] = -11'b00000110100; // -52
storage[3379] = -11'b00000110101; // -53
storage[3380] = -11'b00000100101; // -37
storage[3381] =  11'b00000001110; // 14
storage[3382] = -11'b00001111110; // -126
storage[3383] =  11'b00000001011; // 11
storage[3384] = -11'b00000001111; // -15
storage[3385] = -11'b00000010010; // -18
storage[3386] =  11'b00000000010; // 2
storage[3387] = -11'b00000111011; // -59
storage[3388] =  11'b00000001111; // 15
storage[3389] =  11'b00000000111; // 7
storage[3390] = -11'b00000011001; // -25
storage[3391] = -11'b00000001001; // -9
storage[3392] =  11'b00000000010; // 2
storage[3393] =  11'b00000100101; // 37
storage[3394] = -11'b00000010011; // -19
storage[3395] =  11'b00000110010; // 50
storage[3396] = -11'b00000011100; // -28
storage[3397] =  11'b00001000110; // 70
storage[3398] =  11'b00000100100; // 36
storage[3399] = -11'b00000011101; // -29
storage[3400] =  11'b00001011000; // 88
storage[3401] = -11'b00000100010; // -34
storage[3402] =  11'b00000100011; // 35
storage[3403] =  11'b00000111100; // 60
storage[3404] = -11'b00000101000; // -40
storage[3405] = -11'b00001101101; // -109
storage[3406] =  11'b00000010000; // 16
storage[3407] = -11'b00000011011; // -27
storage[3408] = -11'b00000001010; // -10
storage[3409] = -11'b00000001110; // -14
storage[3410] = -11'b00001011111; // -95
storage[3411] = -11'b00000011001; // -25
storage[3412] = -11'b00000011001; // -25
storage[3413] = -11'b00000000011; // -3
storage[3414] =  11'b00001011100; // 92
storage[3415] =  11'b00000001111; // 15
storage[3416] =  11'b00000011000; // 24
storage[3417] =  11'b00000101101; // 45
storage[3418] = -11'b00000110011; // -51
storage[3419] =  11'b00000111101; // 61
storage[3420] =  11'b00000010101; // 21
storage[3421] = -11'b00000000111; // -7
storage[3422] =  11'b00000010010; // 18
storage[3423] =  11'b00000001011; // 11
storage[3424] =  11'b00001010110; // 86
storage[3425] =  11'b00000010011; // 19
storage[3426] =  11'b00000111100; // 60
storage[3427] = -11'b00000010011; // -19
storage[3428] = -11'b00000110100; // -52
storage[3429] = -11'b00000110111; // -55
storage[3430] = -11'b00000100001; // -33
storage[3431] = -11'b00000000100; // -4
storage[3432] = -11'b00000001100; // -12
storage[3433] =  11'b00000011110; // 30
storage[3434] =  11'b00000010010; // 18
storage[3435] =  11'b00001000111; // 71
storage[3436] = -11'b00000111100; // -60
storage[3437] = -11'b00001000111; // -71
storage[3438] =  11'b00000011100; // 28
storage[3439] = -11'b00001011011; // -91
storage[3440] =  11'b00000011010; // 26
storage[3441] = -11'b00001000010; // -66
storage[3442] =  11'b00000100111; // 39
storage[3443] = -11'b00000001011; // -11
storage[3444] =  11'b00000010100; // 20
storage[3445] =  11'b00001000101; // 69
storage[3446] =  11'b00000010011; // 19
storage[3447] =  11'b00000110000; // 48
storage[3448] = -11'b00000100100; // -36
storage[3449] = -11'b00000001001; // -9
storage[3450] = -11'b00000010111; // -23
storage[3451] =  11'b00000100010; // 34
storage[3452] = -11'b00010000111; // -135
storage[3453] = -11'b00001101110; // -110
storage[3454] = -11'b00010100100; // -164
storage[3455] = -11'b00001001101; // -77
storage[3456] = -11'b00001101001; // -105
storage[3457] =  11'b00000011101; // 29
storage[3458] = -11'b00000001101; // -13
storage[3459] = -11'b00000000101; // -5
storage[3460] =  11'b00000110000; // 48
storage[3461] =  11'b00000000000; // 0
storage[3462] =  11'b00000100001; // 33
storage[3463] =  11'b00000111001; // 57
storage[3464] = -11'b00000000100; // -4
storage[3465] = -11'b00000000001; // -1
storage[3466] = -11'b00001111111; // -127
storage[3467] = -11'b00001000001; // -65
storage[3468] =  11'b00000001001; // 9
storage[3469] = -11'b00000111101; // -61
storage[3470] = -11'b00001010010; // -82
storage[3471] =  11'b00000010000; // 16
storage[3472] = -11'b00001010101; // -85
storage[3473] =  11'b00000101111; // 47
storage[3474] =  11'b00000001100; // 12
storage[3475] = -11'b00000100100; // -36
storage[3476] = -11'b00000000110; // -6
storage[3477] =  11'b00000001101; // 13
storage[3478] =  11'b00001001111; // 79
storage[3479] = -11'b00000011110; // -30
storage[3480] = -11'b00000101010; // -42
storage[3481] =  11'b00001001011; // 75
storage[3482] = -11'b00000010100; // -20
storage[3483] = -11'b00000111001; // -57
storage[3484] = -11'b00000101111; // -47
storage[3485] =  11'b00000000010; // 2
storage[3486] =  11'b00000110011; // 51
storage[3487] =  11'b00000010011; // 19
storage[3488] =  11'b00000101111; // 47
storage[3489] =  11'b00001001011; // 75
storage[3490] =  11'b00000100000; // 32
storage[3491] = -11'b00001011011; // -91
storage[3492] =  11'b00001100010; // 98
storage[3493] =  11'b00000101100; // 44
storage[3494] =  11'b00000101101; // 45
storage[3495] =  11'b00010011110; // 158
storage[3496] = -11'b00000000010; // -2
storage[3497] =  11'b00000000111; // 7
storage[3498] =  11'b00001100011; // 99
storage[3499] = -11'b00000101111; // -47
storage[3500] =  11'b00000000010; // 2
storage[3501] =  11'b00001000001; // 65
storage[3502] =  11'b00000100110; // 38
storage[3503] =  11'b00000101010; // 42
storage[3504] = -11'b00000000100; // -4
storage[3505] = -11'b00000100100; // -36
storage[3506] =  11'b00000110011; // 51
storage[3507] =  11'b00000000001; // 1
storage[3508] = -11'b00000111101; // -61
storage[3509] =  11'b00000110001; // 49
storage[3510] = -11'b00000001100; // -12
storage[3511] =  11'b00000001011; // 11
storage[3512] =  11'b00000011011; // 27
storage[3513] = -11'b00000110010; // -50
storage[3514] =  11'b00000010110; // 22
storage[3515] =  11'b00000000000; // 0
storage[3516] =  11'b00000001010; // 10
storage[3517] = -11'b00000101011; // -43
storage[3518] =  11'b00000001000; // 8
storage[3519] =  11'b00000000100; // 4
storage[3520] =  11'b00000000111; // 7
storage[3521] =  11'b00000000010; // 2
storage[3522] =  11'b00000010110; // 22
storage[3523] =  11'b00001000111; // 71
storage[3524] =  11'b00000001001; // 9
storage[3525] =  11'b00000000001; // 1
storage[3526] =  11'b00000000001; // 1
storage[3527] =  11'b00000010100; // 20
storage[3528] =  11'b00001001001; // 73
storage[3529] = -11'b00001000111; // -71
storage[3530] = -11'b00000010000; // -16
storage[3531] =  11'b00000110111; // 55
storage[3532] = -11'b00000110001; // -49
storage[3533] = -11'b00000010000; // -16
storage[3534] =  11'b00000010110; // 22
storage[3535] =  11'b00000110110; // 54
storage[3536] =  11'b00000010111; // 23
storage[3537] =  11'b00000010011; // 19
storage[3538] =  11'b00001101110; // 110
storage[3539] = -11'b00000001111; // -15
storage[3540] = -11'b00000010001; // -17
storage[3541] = -11'b00000101000; // -40
storage[3542] =  11'b00001100110; // 102
storage[3543] =  11'b00000010000; // 16
storage[3544] =  11'b00000110000; // 48
storage[3545] =  11'b00001010101; // 85
storage[3546] = -11'b00000001110; // -14
storage[3547] =  11'b00000100111; // 39
storage[3548] =  11'b00000001011; // 11
storage[3549] =  11'b00001000011; // 67
storage[3550] = -11'b00000111101; // -61
storage[3551] = -11'b00000011000; // -24
storage[3552] =  11'b00000000111; // 7
storage[3553] =  11'b00000000010; // 2
storage[3554] =  11'b00000111010; // 58
storage[3555] =  11'b00000111000; // 56
storage[3556] = -11'b00000010110; // -22
storage[3557] =  11'b00000110010; // 50
storage[3558] =  11'b00000001000; // 8
storage[3559] =  11'b00000001100; // 12
storage[3560] =  11'b00001000000; // 64
storage[3561] =  11'b00000100011; // 35
storage[3562] = -11'b00000011101; // -29
storage[3563] = -11'b00000100001; // -33
storage[3564] = -11'b00000101010; // -42
storage[3565] = -11'b00000010000; // -16
storage[3566] = -11'b00001100001; // -97
storage[3567] =  11'b00000001010; // 10
storage[3568] = -11'b00000000101; // -5
storage[3569] = -11'b00000110110; // -54
storage[3570] =  11'b00000000011; // 3
storage[3571] =  11'b00000110111; // 55
storage[3572] = -11'b00011001010; // -202
storage[3573] = -11'b00001010001; // -81
storage[3574] = -11'b00001011111; // -95
storage[3575] =  11'b00000001110; // 14
storage[3576] = -11'b00000110010; // -50
storage[3577] = -11'b00010001010; // -138
storage[3578] =  11'b00000010110; // 22
storage[3579] = -11'b00001000111; // -71
storage[3580] =  11'b00000000010; // 2
storage[3581] =  11'b00000010001; // 17
storage[3582] =  11'b00001011100; // 92
storage[3583] = -11'b00001000100; // -68
storage[3584] = -11'b00000001111; // -15
storage[3585] =  11'b00000010111; // 23
storage[3586] = -11'b00001110001; // -113
storage[3587] = -11'b00000011110; // -30
storage[3588] =  11'b00000000011; // 3
storage[3589] =  11'b00000110011; // 51
storage[3590] =  11'b00000010010; // 18
storage[3591] =  11'b00000001011; // 11
storage[3592] = -11'b00001010011; // -83
storage[3593] =  11'b00000011000; // 24
storage[3594] =  11'b00001000000; // 64
storage[3595] = -11'b00001010111; // -87
storage[3596] = -11'b00000001111; // -15
storage[3597] =  11'b00000000111; // 7
storage[3598] = -11'b00010000010; // -130
storage[3599] = -11'b00011110011; // -243
storage[3600] = -11'b00000001011; // -11
storage[3601] =  11'b00000010110; // 22
storage[3602] =  11'b00000110111; // 55
storage[3603] =  11'b00000100001; // 33
storage[3604] = -11'b00000001111; // -15
storage[3605] =  11'b00000000110; // 6
storage[3606] =  11'b00001001111; // 79
storage[3607] = -11'b00001110110; // -118
storage[3608] = -11'b00000101010; // -42
storage[3609] =  11'b00000100101; // 37
storage[3610] = -11'b00000111010; // -58
storage[3611] =  11'b00001000001; // 65
storage[3612] =  11'b00000100010; // 34
storage[3613] =  11'b00001000101; // 69
storage[3614] =  11'b00001001000; // 72
storage[3615] = -11'b00000001110; // -14
storage[3616] = -11'b00000011010; // -26
storage[3617] = -11'b00000000001; // -1
storage[3618] =  11'b00000011101; // 29
storage[3619] =  11'b00001101100; // 108
storage[3620] = -11'b00001011101; // -93
storage[3621] = -11'b00000111001; // -57
storage[3622] =  11'b00000110111; // 55
storage[3623] = -11'b00000000100; // -4
storage[3624] =  11'b00000001010; // 10
storage[3625] = -11'b00000100101; // -37
storage[3626] =  11'b00001000010; // 66
storage[3627] = -11'b00000010011; // -19
storage[3628] = -11'b00000111110; // -62
storage[3629] = -11'b00000100010; // -34
storage[3630] =  11'b00000101000; // 40
storage[3631] = -11'b00000001011; // -11
storage[3632] =  11'b00000001000; // 8
storage[3633] = -11'b00000101000; // -40
storage[3634] = -11'b00000111010; // -58
storage[3635] =  11'b00000000001; // 1
storage[3636] =  11'b00000000000; // 0
storage[3637] = -11'b00000001101; // -13
storage[3638] = -11'b00000010011; // -19
storage[3639] =  11'b00000010011; // 19
storage[3640] = -11'b00000000010; // -2
storage[3641] =  11'b00000001101; // 13
storage[3642] =  11'b00000001001; // 9
storage[3643] =  11'b00000101100; // 44
storage[3644] =  11'b00000010001; // 17
storage[3645] = -11'b00000011001; // -25
storage[3646] = -11'b00001011011; // -91
storage[3647] =  11'b00000000000; // 0
storage[3648] = -11'b00000000110; // -6
storage[3649] = -11'b00010000000; // -128
storage[3650] =  11'b00000011010; // 26
storage[3651] =  11'b00000010010; // 18
storage[3652] = -11'b00001010100; // -84
storage[3653] = -11'b00000011000; // -24
storage[3654] = -11'b00010100110; // -166
storage[3655] = -11'b00001011000; // -88
storage[3656] = -11'b00000101100; // -44
storage[3657] =  11'b00000000011; // 3
storage[3658] = -11'b00000001010; // -10
storage[3659] = -11'b00001010111; // -87
storage[3660] =  11'b00000001001; // 9
storage[3661] = -11'b00001101000; // -104
storage[3662] = -11'b00010011100; // -156
storage[3663] = -11'b00001011010; // -90
storage[3664] =  11'b00000011101; // 29
storage[3665] =  11'b00000110001; // 49
storage[3666] =  11'b00000001010; // 10
storage[3667] =  11'b00000000001; // 1
storage[3668] =  11'b00000011101; // 29
storage[3669] = -11'b00000101001; // -41
storage[3670] =  11'b00000101011; // 43
storage[3671] =  11'b00000101111; // 47
storage[3672] = -11'b00000010110; // -22
storage[3673] = -11'b00000011001; // -25
storage[3674] = -11'b00001110010; // -114
storage[3675] =  11'b00000000110; // 6
storage[3676] = -11'b00000001010; // -10
storage[3677] = -11'b00000111111; // -63
storage[3678] =  11'b00000001001; // 9
storage[3679] =  11'b00000010100; // 20
storage[3680] =  11'b00000100001; // 33
storage[3681] =  11'b00000000011; // 3
storage[3682] = -11'b00010010101; // -149
storage[3683] = -11'b00001000011; // -67
storage[3684] =  11'b00000100110; // 38
storage[3685] = -11'b00000110001; // -49
storage[3686] = -11'b00000110000; // -48
storage[3687] =  11'b00000101000; // 40
storage[3688] = -11'b00000000100; // -4
storage[3689] = -11'b00000100110; // -38
storage[3690] =  11'b00000001011; // 11
storage[3691] =  11'b00001011000; // 88
storage[3692] =  11'b00000011101; // 29
storage[3693] =  11'b00000011101; // 29
storage[3694] =  11'b00000110000; // 48
storage[3695] =  11'b00000011101; // 29
storage[3696] =  11'b00000000011; // 3
storage[3697] = -11'b00000110010; // -50
storage[3698] = -11'b00000110111; // -55
storage[3699] = -11'b00000000011; // -3
storage[3700] =  11'b00000000110; // 6
storage[3701] = -11'b00000001111; // -15
storage[3702] = -11'b00000011000; // -24
storage[3703] =  11'b00000100001; // 33
storage[3704] =  11'b00000010001; // 17
storage[3705] = -11'b00001001000; // -72
storage[3706] =  11'b00000001001; // 9
storage[3707] = -11'b00000011100; // -28
storage[3708] = -11'b00001110010; // -114
storage[3709] = -11'b00000111010; // -58
storage[3710] = -11'b00000010011; // -19
storage[3711] =  11'b00000100010; // 34
storage[3712] =  11'b00000010010; // 18
storage[3713] = -11'b00000011000; // -24
storage[3714] = -11'b00001010101; // -85
storage[3715] =  11'b00001011011; // 91
storage[3716] =  11'b00000111010; // 58
storage[3717] = -11'b00000000100; // -4
storage[3718] = -11'b00001001101; // -77
storage[3719] =  11'b00000001000; // 8
storage[3720] = -11'b00001000101; // -69
storage[3721] =  11'b00001000111; // 71
storage[3722] =  11'b00000001110; // 14
storage[3723] = -11'b00010010100; // -148
storage[3724] =  11'b00001010101; // 85
storage[3725] =  11'b00000111101; // 61
storage[3726] = -11'b00000010010; // -18
storage[3727] =  11'b00000010110; // 22
storage[3728] =  11'b00000101110; // 46
storage[3729] = -11'b00000001001; // -9
storage[3730] =  11'b00000001100; // 12
storage[3731] =  11'b00001000101; // 69
storage[3732] = -11'b00000010110; // -22
storage[3733] = -11'b00000010010; // -18
storage[3734] =  11'b00001001001; // 73
storage[3735] = -11'b00000001001; // -9
storage[3736] = -11'b00000111100; // -60
storage[3737] = -11'b00000110010; // -50
storage[3738] =  11'b00000110100; // 52
storage[3739] = -11'b00000111110; // -62
storage[3740] =  11'b00000001011; // 11
storage[3741] =  11'b00001011111; // 95
storage[3742] = -11'b00000111000; // -56
storage[3743] =  11'b00001000011; // 67
storage[3744] =  11'b00000110110; // 54
storage[3745] = -11'b00000000010; // -2
storage[3746] =  11'b00001000101; // 69
storage[3747] =  11'b00000000111; // 7
storage[3748] =  11'b00000011111; // 31
storage[3749] =  11'b00000101110; // 46
storage[3750] = -11'b00000000111; // -7
storage[3751] = -11'b00000100100; // -36
storage[3752] = -11'b00000001011; // -11
storage[3753] = -11'b00000100111; // -39
storage[3754] =  11'b00000011110; // 30
storage[3755] = -11'b00000010101; // -21
storage[3756] = -11'b00000111010; // -58
storage[3757] =  11'b00000000110; // 6
storage[3758] = -11'b00000001011; // -11
storage[3759] = -11'b00000100100; // -36
storage[3760] =  11'b00000010111; // 23
storage[3761] =  11'b00000001100; // 12
storage[3762] = -11'b00000011001; // -25
storage[3763] = -11'b00001011010; // -90
storage[3764] = -11'b00000011101; // -29
storage[3765] =  11'b00000001000; // 8
storage[3766] = -11'b00001100110; // -102
storage[3767] =  11'b00000001111; // 15
storage[3768] =  11'b00000000110; // 6
storage[3769] = -11'b00000011100; // -28
storage[3770] = -11'b00011100100; // -228
storage[3771] =  11'b00000100011; // 35
storage[3772] =  11'b00000110001; // 49
storage[3773] =  11'b00001110111; // 119
storage[3774] =  11'b00001010001; // 81
storage[3775] = -11'b00001001100; // -76
storage[3776] =  11'b00000011000; // 24
storage[3777] = -11'b00000001010; // -10
storage[3778] = -11'b00000011011; // -27
storage[3779] = -11'b00000101000; // -40
storage[3780] = -11'b00000100101; // -37
storage[3781] = -11'b00000100101; // -37
storage[3782] = -11'b00010001101; // -141
storage[3783] = -11'b00000011011; // -27
storage[3784] = -11'b00010000001; // -129
storage[3785] = -11'b00000010111; // -23
storage[3786] =  11'b00000110100; // 52
storage[3787] =  11'b00000010000; // 16
storage[3788] =  11'b00000000001; // 1
storage[3789] = -11'b00000110110; // -54
storage[3790] = -11'b00000101110; // -46
storage[3791] =  11'b00000010001; // 17
storage[3792] =  11'b00000000010; // 2
storage[3793] = -11'b00001100100; // -100
storage[3794] = -11'b00000110011; // -51
storage[3795] =  11'b00001000111; // 71
storage[3796] = -11'b00000000011; // -3
storage[3797] =  11'b00000011010; // 26
storage[3798] =  11'b00000000010; // 2
storage[3799] = -11'b00010010100; // -148
storage[3800] = -11'b00001001011; // -75
storage[3801] =  11'b00001000001; // 65
storage[3802] = -11'b00010010110; // -150
storage[3803] = -11'b00000101000; // -40
storage[3804] =  11'b00001001000; // 72
storage[3805] =  11'b00000000101; // 5
storage[3806] = -11'b00001111110; // -126
storage[3807] =  11'b00000001101; // 13
storage[3808] = -11'b00010100001; // -161
storage[3809] = -11'b00000010001; // -17
storage[3810] =  11'b00000111010; // 58
storage[3811] = -11'b00000000001; // -1
storage[3812] =  11'b00000011101; // 29
storage[3813] =  11'b00000101010; // 42
storage[3814] =  11'b00001001010; // 74
storage[3815] = -11'b00000011010; // -26
storage[3816] = -11'b00000011000; // -24
storage[3817] = -11'b00000001011; // -11
storage[3818] =  11'b00000010001; // 17
storage[3819] =  11'b00001000111; // 71
storage[3820] = -11'b00000100111; // -39
storage[3821] = -11'b00000100100; // -36
storage[3822] =  11'b00000001111; // 15
storage[3823] = -11'b00001111100; // -124
storage[3824] = -11'b00000011001; // -25
storage[3825] = -11'b00000010001; // -17
storage[3826] =  11'b00001011011; // 91
storage[3827] =  11'b00000101000; // 40
storage[3828] =  11'b00000001110; // 14
storage[3829] = -11'b00000011011; // -27
storage[3830] =  11'b00000011001; // 25
storage[3831] = -11'b00000101100; // -44
storage[3832] = -11'b00001100100; // -100
storage[3833] = -11'b00000111111; // -63
storage[3834] = -11'b00000011001; // -25
storage[3835] =  11'b00000100010; // 34
storage[3836] =  11'b00000011110; // 30
storage[3837] =  11'b00001011100; // 92
storage[3838] = -11'b00000100011; // -35
storage[3839] =  11'b00000010001; // 17
storage[3840] =  11'b00000011100; // 28
storage[3841] = -11'b00000001010; // -10
storage[3842] =  11'b00000001110; // 14
storage[3843] =  11'b00000011001; // 25
storage[3844] = -11'b00000010000; // -16
storage[3845] = -11'b00001011000; // -88
storage[3846] = -11'b00000010101; // -21
storage[3847] = -11'b00000010100; // -20
storage[3848] =  11'b00000100110; // 38
storage[3849] =  11'b00000101010; // 42
storage[3850] = -11'b00000011001; // -25
storage[3851] = -11'b00000000100; // -4
storage[3852] =  11'b00000111101; // 61
storage[3853] =  11'b00000001001; // 9
storage[3854] =  11'b00000101000; // 40
storage[3855] =  11'b00000000100; // 4
storage[3856] = -11'b00000110111; // -55
storage[3857] = -11'b00000010000; // -16
storage[3858] =  11'b00000011101; // 29
storage[3859] =  11'b00000100000; // 32
storage[3860] =  11'b00000110011; // 51
storage[3861] =  11'b00001100001; // 97
storage[3862] =  11'b00000100101; // 37
storage[3863] =  11'b00001010010; // 82
storage[3864] =  11'b00000011111; // 31
storage[3865] = -11'b00000010110; // -22
storage[3866] =  11'b00000010010; // 18
storage[3867] =  11'b00000011000; // 24
storage[3868] =  11'b00000001110; // 14
storage[3869] =  11'b00001010000; // 80
storage[3870] =  11'b00000100011; // 35
storage[3871] = -11'b00001000010; // -66
storage[3872] =  11'b00000110110; // 54
storage[3873] =  11'b00000000010; // 2
storage[3874] = -11'b00000010010; // -18
storage[3875] =  11'b00000010101; // 21
storage[3876] =  11'b00000101111; // 47
storage[3877] = -11'b00001010000; // -80
storage[3878] = -11'b00000010011; // -19
storage[3879] =  11'b00000001101; // 13
storage[3880] =  11'b00000101100; // 44
storage[3881] =  11'b00000011011; // 27
storage[3882] =  11'b00001000111; // 71
storage[3883] =  11'b00000100111; // 39
storage[3884] =  11'b00000001110; // 14
storage[3885] =  11'b00000101011; // 43
storage[3886] =  11'b00001000001; // 65
storage[3887] =  11'b00000101010; // 42
storage[3888] = -11'b00000001101; // -13
storage[3889] = -11'b00001001111; // -79
storage[3890] =  11'b00000000100; // 4
storage[3891] =  11'b00000110010; // 50
storage[3892] = -11'b00000001011; // -11
storage[3893] =  11'b00000001100; // 12
storage[3894] =  11'b00000000101; // 5
storage[3895] = -11'b00000101000; // -40
storage[3896] = -11'b00000110101; // -53
storage[3897] = -11'b00000001010; // -10
storage[3898] = -11'b00010000100; // -132
storage[3899] = -11'b00000000001; // -1
storage[3900] =  11'b00000100010; // 34
storage[3901] = -11'b00001001000; // -72
storage[3902] = -11'b00000000010; // -2
storage[3903] =  11'b00000111000; // 56
storage[3904] = -11'b00000011000; // -24
storage[3905] =  11'b00000010101; // 21
storage[3906] =  11'b00000011010; // 26
storage[3907] = -11'b00000100101; // -37
storage[3908] =  11'b00000001101; // 13
storage[3909] = -11'b00010010001; // -145
storage[3910] = -11'b00000010010; // -18
storage[3911] = -11'b00001110011; // -115
storage[3912] = -11'b00000110010; // -50
storage[3913] =  11'b00000101010; // 42
storage[3914] = -11'b00000101111; // -47
storage[3915] = -11'b00001010111; // -87
storage[3916] = -11'b00000101001; // -41
storage[3917] = -11'b00001001111; // -79
storage[3918] = -11'b00000010010; // -18
storage[3919] =  11'b00000000110; // 6
storage[3920] =  11'b00000010010; // 18
storage[3921] = -11'b00000000100; // -4
storage[3922] = -11'b00000001001; // -9
storage[3923] =  11'b00000010000; // 16
storage[3924] = -11'b00000101011; // -43
storage[3925] =  11'b00001001100; // 76
storage[3926] =  11'b00000011011; // 27
storage[3927] =  11'b00000110010; // 50
storage[3928] =  11'b00000000111; // 7
storage[3929] = -11'b00000000110; // -6
storage[3930] = -11'b00000011110; // -30
storage[3931] =  11'b00000011100; // 28
storage[3932] = -11'b00000000011; // -3
storage[3933] = -11'b00000010101; // -21
storage[3934] = -11'b00000101011; // -43
storage[3935] = -11'b00000001000; // -8
storage[3936] =  11'b00000101011; // 43
storage[3937] = -11'b00001101001; // -105
storage[3938] = -11'b00000101100; // -44
storage[3939] = -11'b00000111110; // -62
storage[3940] = -11'b00000101100; // -44
storage[3941] = -11'b00000011111; // -31
storage[3942] = -11'b00000110110; // -54
storage[3943] = -11'b00000001011; // -11
storage[3944] = -11'b00000001101; // -13
storage[3945] =  11'b00000001001; // 9
storage[3946] = -11'b00000001011; // -11
storage[3947] = -11'b00000001101; // -13
storage[3948] = -11'b00001011010; // -90
storage[3949] =  11'b00000000001; // 1
storage[3950] =  11'b00000001001; // 9
storage[3951] = -11'b00000010100; // -20
storage[3952] = -11'b00000001101; // -13
storage[3953] = -11'b00000010001; // -17
storage[3954] =  11'b00000010001; // 17
storage[3955] =  11'b00000110100; // 52
storage[3956] = -11'b00000010000; // -16
storage[3957] = -11'b00001111000; // -120
storage[3958] =  11'b00000001101; // 13
storage[3959] =  11'b00000100001; // 33
storage[3960] = -11'b00000011100; // -28
storage[3961] =  11'b00000011100; // 28
storage[3962] = -11'b00000100101; // -37
storage[3963] = -11'b00000010011; // -19
storage[3964] =  11'b00001000000; // 64
storage[3965] =  11'b00000000011; // 3
storage[3966] = -11'b00000010000; // -16
storage[3967] =  11'b00000111001; // 57
storage[3968] =  11'b00000011011; // 27
storage[3969] = -11'b00000101101; // -45
storage[3970] = -11'b00001000110; // -70
storage[3971] =  11'b00000000111; // 7
storage[3972] =  11'b00000110000; // 48
storage[3973] = -11'b00000001111; // -15
storage[3974] =  11'b00000000010; // 2
storage[3975] =  11'b00000001010; // 10
storage[3976] =  11'b00000001101; // 13
storage[3977] =  11'b00000110101; // 53
storage[3978] = -11'b00000101110; // -46
storage[3979] = -11'b00000011110; // -30
storage[3980] = -11'b00000010110; // -22
storage[3981] =  11'b00000001100; // 12
storage[3982] =  11'b00000000110; // 6
storage[3983] = -11'b00000100010; // -34
storage[3984] = -11'b00000001101; // -13
storage[3985] = -11'b00000011111; // -31
storage[3986] =  11'b00000001011; // 11
storage[3987] = -11'b00000000100; // -4
storage[3988] = -11'b00000011011; // -27
storage[3989] =  11'b00000011001; // 25
storage[3990] = -11'b00001000000; // -64
storage[3991] = -11'b00000000001; // -1
storage[3992] =  11'b00000000110; // 6
storage[3993] =  11'b00000100101; // 37
storage[3994] =  11'b00000000101; // 5
storage[3995] = -11'b00000001110; // -14
storage[3996] =  11'b00000001110; // 14
storage[3997] =  11'b00000101011; // 43
storage[3998] = -11'b00000100010; // -34
storage[3999] = -11'b00000011000; // -24
storage[4000] = -11'b00001110111; // -119
storage[4001] = -11'b00001011111; // -95
storage[4002] =  11'b00000011111; // 31
storage[4003] = -11'b00000110101; // -53
storage[4004] = -11'b00000001000; // -8
storage[4005] =  11'b00001000001; // 65
storage[4006] = -11'b00000110101; // -53
storage[4007] = -11'b00000000001; // -1
storage[4008] =  11'b00000110010; // 50
storage[4009] =  11'b00000000000; // 0
storage[4010] =  11'b00000010101; // 21
storage[4011] = -11'b00000001001; // -9
storage[4012] =  11'b00000111111; // 63
storage[4013] =  11'b00000010101; // 21
storage[4014] = -11'b00000011011; // -27
storage[4015] = -11'b00000010101; // -21
storage[4016] = -11'b00001101101; // -109
storage[4017] = -11'b00000101000; // -40
storage[4018] = -11'b00000000110; // -6
storage[4019] = -11'b00000110011; // -51
storage[4020] = -11'b00000000100; // -4
storage[4021] =  11'b00000010001; // 17
storage[4022] =  11'b00000111011; // 59
storage[4023] =  11'b00000101100; // 44
storage[4024] =  11'b00000011011; // 27
storage[4025] =  11'b00000100111; // 39
storage[4026] =  11'b00000011111; // 31
storage[4027] = -11'b00000000101; // -5
storage[4028] =  11'b00000111101; // 61
storage[4029] =  11'b00000000101; // 5
storage[4030] = -11'b00000001111; // -15
storage[4031] =  11'b00000010101; // 21
storage[4032] = -11'b00010010010; // -146
storage[4033] =  11'b00000000011; // 3
storage[4034] =  11'b00000101100; // 44
storage[4035] = -11'b00000001010; // -10
storage[4036] = -11'b00000000111; // -7
storage[4037] =  11'b00000110110; // 54
storage[4038] =  11'b00000101101; // 45
storage[4039] =  11'b00000100101; // 37
storage[4040] =  11'b00000111001; // 57
storage[4041] =  11'b00000001100; // 12
storage[4042] = -11'b00000101000; // -40
storage[4043] = -11'b00000111110; // -62
storage[4044] =  11'b00000000100; // 4
storage[4045] =  11'b00001110100; // 116
storage[4046] =  11'b00000000001; // 1
storage[4047] =  11'b00000001000; // 8
storage[4048] =  11'b00001001100; // 76
storage[4049] =  11'b00000010111; // 23
storage[4050] = -11'b00000000010; // -2
storage[4051] =  11'b00001010101; // 85
storage[4052] = -11'b00000110100; // -52
storage[4053] =  11'b00000011011; // 27
storage[4054] = -11'b00001010010; // -82
storage[4055] = -11'b00001001110; // -78
storage[4056] =  11'b00001000100; // 68
storage[4057] = -11'b00000001011; // -11
storage[4058] = -11'b00001001111; // -79
storage[4059] = -11'b00000110101; // -53
storage[4060] = -11'b00010000100; // -132
storage[4061] = -11'b00001100111; // -103
storage[4062] = -11'b00000011110; // -30
storage[4063] = -11'b00010010011; // -147
storage[4064] = -11'b00000100010; // -34
storage[4065] =  11'b00000011110; // 30
storage[4066] = -11'b00000111101; // -61
storage[4067] = -11'b00000101110; // -46
storage[4068] = -11'b00000100111; // -39
storage[4069] =  11'b00000100001; // 33
storage[4070] =  11'b00000001101; // 13
storage[4071] =  11'b00000000101; // 5
storage[4072] =  11'b00000110001; // 49
storage[4073] =  11'b00000000000; // 0
storage[4074] = -11'b00000011100; // -28
storage[4075] = -11'b00000110011; // -51
storage[4076] = -11'b00000101111; // -47
storage[4077] = -11'b00000010110; // -22
storage[4078] =  11'b00000001011; // 11
storage[4079] = -11'b00001001100; // -76
storage[4080] =  11'b00000011010; // 26
storage[4081] = -11'b00000111100; // -60
storage[4082] = -11'b00000010101; // -21
storage[4083] =  11'b00000100000; // 32
storage[4084] = -11'b00000010110; // -22
storage[4085] =  11'b00001010110; // 86
storage[4086] = -11'b00000101001; // -41
storage[4087] =  11'b00000010101; // 21
storage[4088] =  11'b00000011100; // 28
storage[4089] = -11'b00000101111; // -47
storage[4090] = -11'b00000010011; // -19
storage[4091] = -11'b00000101100; // -44
storage[4092] = -11'b00000101010; // -42
storage[4093] = -11'b00001101010; // -106
storage[4094] = -11'b00000111100; // -60
storage[4095] =  11'b00000001100; // 12
storage[4096] =  11'b00000000100; // 4
storage[4097] = -11'b00000000010; // -2
storage[4098] =  11'b00000100000; // 32
storage[4099] = -11'b00000010010; // -18
storage[4100] = -11'b00000010000; // -16
storage[4101] =  11'b00000111000; // 56
storage[4102] = -11'b00000010111; // -23
storage[4103] =  11'b00000011011; // 27
storage[4104] =  11'b00001000101; // 69
storage[4105] = -11'b00000001000; // -8
storage[4106] =  11'b00000110101; // 53
storage[4107] =  11'b00000000000; // 0
storage[4108] = -11'b00000001010; // -10
storage[4109] =  11'b00000001111; // 15
storage[4110] =  11'b00000011011; // 27
storage[4111] = -11'b00001100111; // -103
storage[4112] = -11'b00000110101; // -53
storage[4113] = -11'b00000100111; // -39
storage[4114] = -11'b00000000111; // -7
storage[4115] = -11'b00000111010; // -58
storage[4116] = -11'b00000011001; // -25
storage[4117] = -11'b00000010100; // -20
storage[4118] =  11'b00000100110; // 38
storage[4119] = -11'b00000010110; // -22
storage[4120] = -11'b00001110011; // -115
storage[4121] = -11'b00001011001; // -89
storage[4122] =  11'b00000010001; // 17
storage[4123] = -11'b00000000111; // -7
storage[4124] = -11'b00000011110; // -30
storage[4125] = -11'b00000110111; // -55
storage[4126] =  11'b00001000100; // 68
storage[4127] =  11'b00001010101; // 85
storage[4128] =  11'b00000011001; // 25
storage[4129] =  11'b00001000110; // 70
storage[4130] =  11'b00000011001; // 25
storage[4131] = -11'b00000010111; // -23
storage[4132] =  11'b00000000000; // 0
storage[4133] =  11'b00000001110; // 14
storage[4134] =  11'b00000101100; // 44
storage[4135] =  11'b00000001000; // 8
storage[4136] = -11'b00000001001; // -9
storage[4137] = -11'b00000001001; // -9
storage[4138] =  11'b00000011011; // 27
storage[4139] =  11'b00000111101; // 61
storage[4140] = -11'b00000000101; // -5
storage[4141] = -11'b00000000001; // -1
storage[4142] = -11'b00000010011; // -19
storage[4143] = -11'b00000001110; // -14
storage[4144] =  11'b00000010001; // 17
storage[4145] =  11'b00000000101; // 5
storage[4146] =  11'b00000010101; // 21
storage[4147] =  11'b00000001000; // 8
storage[4148] =  11'b00000011110; // 30
storage[4149] = -11'b00010001110; // -142
storage[4150] =  11'b00000110110; // 54
storage[4151] =  11'b00000011000; // 24
storage[4152] = -11'b00000111000; // -56
storage[4153] = -11'b00000100100; // -36
storage[4154] =  11'b00000100110; // 38
storage[4155] = -11'b00001100010; // -98
storage[4156] = -11'b00000000111; // -7
storage[4157] = -11'b00000000001; // -1
storage[4158] = -11'b00000101011; // -43
storage[4159] =  11'b00000001011; // 11
storage[4160] =  11'b00000101010; // 42
storage[4161] =  11'b00000010000; // 16
storage[4162] =  11'b00000001100; // 12
storage[4163] =  11'b00000101000; // 40
storage[4164] =  11'b00000101001; // 41
storage[4165] = -11'b00000000111; // -7
storage[4166] = -11'b00000001000; // -8
storage[4167] = -11'b00000001001; // -9
storage[4168] = -11'b00000101101; // -45
storage[4169] =  11'b00000011010; // 26
storage[4170] = -11'b00000100101; // -37
storage[4171] = -11'b00000101111; // -47
storage[4172] = -11'b00000101111; // -47
storage[4173] = -11'b00001001101; // -77
storage[4174] =  11'b00000111100; // 60
storage[4175] = -11'b00010101000; // -168
storage[4176] = -11'b00001000110; // -70
storage[4177] =  11'b00000000100; // 4
storage[4178] =  11'b00001100001; // 97
storage[4179] = -11'b00000011100; // -28
storage[4180] = -11'b00000000011; // -3
storage[4181] =  11'b00000111001; // 57
storage[4182] =  11'b00000010011; // 19
storage[4183] =  11'b00000110111; // 55
storage[4184] = -11'b00000001101; // -13
storage[4185] = -11'b00000010011; // -19
storage[4186] =  11'b00000110011; // 51
storage[4187] =  11'b00000110111; // 55
storage[4188] = -11'b00000010101; // -21
storage[4189] =  11'b00000100101; // 37
storage[4190] = -11'b00000011000; // -24
storage[4191] = -11'b00000100010; // -34
storage[4192] =  11'b00000011110; // 30
storage[4193] = -11'b00000100011; // -35
storage[4194] = -11'b00000000110; // -6
storage[4195] =  11'b00000010101; // 21
storage[4196] =  11'b00000000010; // 2
storage[4197] =  11'b00000000001; // 1
storage[4198] =  11'b00000001000; // 8
storage[4199] =  11'b00000010110; // 22
storage[4200] =  11'b00000011000; // 24
storage[4201] = -11'b00000100110; // -38
storage[4202] =  11'b00000000000; // 0
storage[4203] =  11'b00000110000; // 48
storage[4204] =  11'b00000000011; // 3
storage[4205] = -11'b00000001010; // -10
storage[4206] =  11'b00001001010; // 74
storage[4207] =  11'b00000000110; // 6
storage[4208] =  11'b00000110110; // 54
storage[4209] =  11'b00000101000; // 40
storage[4210] = -11'b00000010000; // -16
storage[4211] =  11'b00001001101; // 77
storage[4212] =  11'b00000100100; // 36
storage[4213] = -11'b00000110010; // -50
storage[4214] = -11'b00000001000; // -8
storage[4215] = -11'b00000110011; // -51
storage[4216] = -11'b00000001010; // -10
storage[4217] = -11'b00001000111; // -71
storage[4218] = -11'b00000011100; // -28
storage[4219] = -11'b00000000110; // -6
storage[4220] =  11'b00001001101; // 77
storage[4221] = -11'b00000110110; // -54
storage[4222] =  11'b00000011010; // 26
storage[4223] =  11'b00000110000; // 48
storage[4224] = -11'b00000100110; // -38
storage[4225] =  11'b00000011100; // 28
storage[4226] = -11'b00000010110; // -22
storage[4227] =  11'b00000000101; // 5
storage[4228] = -11'b00000011111; // -31
storage[4229] = -11'b00000110101; // -53
storage[4230] = -11'b00000000100; // -4
storage[4231] = -11'b00000111011; // -59
storage[4232] = -11'b00001100000; // -96
storage[4233] = -11'b00010110100; // -180
storage[4234] =  11'b00000001110; // 14
storage[4235] =  11'b00000101010; // 42
storage[4236] =  11'b00000101001; // 41
storage[4237] =  11'b00000001100; // 12
storage[4238] =  11'b00000101001; // 41
storage[4239] =  11'b00000111010; // 58
storage[4240] = -11'b00001101001; // -105
storage[4241] = -11'b00001010111; // -87
storage[4242] = -11'b00001101011; // -107
storage[4243] = -11'b00000011011; // -27
storage[4244] =  11'b00000101001; // 41
storage[4245] =  11'b00000011001; // 25
storage[4246] = -11'b00000100011; // -35
storage[4247] =  11'b00001100100; // 100
storage[4248] =  11'b00001011100; // 92
storage[4249] = -11'b00000110000; // -48
storage[4250] = -11'b00001100001; // -97
storage[4251] =  11'b00000000100; // 4
storage[4252] =  11'b00000110100; // 52
storage[4253] =  11'b00000110000; // 48
storage[4254] = -11'b00000101001; // -41
storage[4255] =  11'b00000011111; // 31
storage[4256] =  11'b00000111101; // 61
storage[4257] =  11'b00000010110; // 22
storage[4258] =  11'b00000110110; // 54
storage[4259] =  11'b00000001100; // 12
storage[4260] =  11'b00000001011; // 11
storage[4261] = -11'b00001000111; // -71
storage[4262] = -11'b00000001110; // -14
storage[4263] = -11'b00000000010; // -2
storage[4264] =  11'b00000001111; // 15
storage[4265] =  11'b00000001110; // 14
storage[4266] = -11'b00100011000; // -280
storage[4267] =  11'b00000011110; // 30
storage[4268] = -11'b00001001100; // -76
storage[4269] = -11'b00001011011; // -91
storage[4270] =  11'b00000101000; // 40
storage[4271] =  11'b00000110100; // 52
storage[4272] =  11'b00000001101; // 13
storage[4273] = -11'b00000010100; // -20
storage[4274] = -11'b00000000001; // -1
storage[4275] =  11'b00000111011; // 59
storage[4276] =  11'b00000000001; // 1
storage[4277] =  11'b00000001010; // 10
storage[4278] =  11'b00001001010; // 74
storage[4279] =  11'b00000000010; // 2
storage[4280] =  11'b00000000000; // 0
storage[4281] = -11'b00000000111; // -7
storage[4282] = -11'b00000010011; // -19
storage[4283] =  11'b00000001111; // 15
storage[4284] =  11'b00001101010; // 106
storage[4285] =  11'b00000100010; // 34
storage[4286] = -11'b00000111110; // -62
storage[4287] = -11'b00010000100; // -132
storage[4288] =  11'b00000000110; // 6
storage[4289] = -11'b00000100111; // -39
storage[4290] = -11'b00010001010; // -138
storage[4291] = -11'b00001111111; // -127
storage[4292] =  11'b00000101101; // 45
storage[4293] = -11'b00000000111; // -7
storage[4294] =  11'b00000000000; // 0
storage[4295] =  11'b00000100101; // 37
storage[4296] =  11'b00000001101; // 13
storage[4297] =  11'b00000001010; // 10
storage[4298] =  11'b00000010101; // 21
storage[4299] =  11'b00000010000; // 16
storage[4300] = -11'b00001100010; // -98
storage[4301] = -11'b00001101110; // -110
storage[4302] =  11'b00001101100; // 108
storage[4303] =  11'b00000011101; // 29
storage[4304] =  11'b00000101111; // 47
storage[4305] = -11'b00000100110; // -38
storage[4306] =  11'b00000011001; // 25
storage[4307] = -11'b00000100011; // -35
storage[4308] = -11'b00000101000; // -40
storage[4309] =  11'b00000011000; // 24
storage[4310] =  11'b00000101110; // 46
storage[4311] =  11'b00000001101; // 13
storage[4312] =  11'b00000110000; // 48
storage[4313] = -11'b00001000110; // -70
storage[4314] = -11'b00000110101; // -53
storage[4315] = -11'b00000010111; // -23
storage[4316] = -11'b00000010100; // -20
storage[4317] = -11'b00000011101; // -29
storage[4318] =  11'b00000011010; // 26
storage[4319] =  11'b00000001010; // 10
storage[4320] = -11'b00000110000; // -48
storage[4321] =  11'b00000001111; // 15
storage[4322] =  11'b00000101101; // 45
storage[4323] =  11'b00000101100; // 44
storage[4324] =  11'b00001000010; // 66
storage[4325] =  11'b00000001000; // 8
storage[4326] =  11'b00000100000; // 32
storage[4327] =  11'b00000010111; // 23
storage[4328] =  11'b00000010001; // 17
storage[4329] = -11'b00000001101; // -13
storage[4330] =  11'b00001001001; // 73
storage[4331] = -11'b00000000110; // -6
storage[4332] =  11'b00000010100; // 20
storage[4333] =  11'b00000110000; // 48
storage[4334] =  11'b00000011000; // 24
storage[4335] = -11'b00000100000; // -32
storage[4336] =  11'b00000010100; // 20
storage[4337] = -11'b00000000010; // -2
storage[4338] = -11'b00000001001; // -9
storage[4339] = -11'b00001101111; // -111
storage[4340] = -11'b00000011000; // -24
storage[4341] =  11'b00000000101; // 5
storage[4342] =  11'b00000000011; // 3
storage[4343] = -11'b00001001000; // -72
storage[4344] =  11'b00000000001; // 1
storage[4345] = -11'b00001000010; // -66
storage[4346] = -11'b00000110100; // -52
storage[4347] = -11'b00000010011; // -19
storage[4348] =  11'b00000000010; // 2
storage[4349] =  11'b00000111111; // 63
storage[4350] =  11'b00000011110; // 30
storage[4351] = -11'b00000001100; // -12
storage[4352] =  11'b00000011110; // 30
storage[4353] = -11'b00000000011; // -3
storage[4354] =  11'b00000101010; // 42
storage[4355] =  11'b00000010011; // 19
storage[4356] =  11'b00000001100; // 12
storage[4357] = -11'b00000010010; // -18
storage[4358] =  11'b00000000011; // 3
storage[4359] =  11'b00000010011; // 19
storage[4360] = -11'b00000010010; // -18
storage[4361] = -11'b00000010111; // -23
storage[4362] = -11'b00000110100; // -52
storage[4363] =  11'b00000010110; // 22
storage[4364] =  11'b00000011111; // 31
storage[4365] =  11'b00001010000; // 80
storage[4366] =  11'b00000010010; // 18
storage[4367] =  11'b00000001000; // 8
storage[4368] =  11'b00000100011; // 35
storage[4369] =  11'b00000100101; // 37
storage[4370] =  11'b00001001111; // 79
storage[4371] =  11'b00000101100; // 44
storage[4372] =  11'b00000110010; // 50
storage[4373] = -11'b00000011010; // -26
storage[4374] =  11'b00000001000; // 8
storage[4375] = -11'b00000010010; // -18
storage[4376] = -11'b00000010100; // -20
storage[4377] = -11'b00000100001; // -33
storage[4378] = -11'b00000011011; // -27
storage[4379] = -11'b00000010100; // -20
storage[4380] = -11'b00000010001; // -17
storage[4381] =  11'b00000011011; // 27
storage[4382] =  11'b00000110000; // 48
storage[4383] =  11'b00000100110; // 38
storage[4384] =  11'b00000000110; // 6
storage[4385] = -11'b00000001000; // -8
storage[4386] =  11'b00000100010; // 34
storage[4387] =  11'b00000100011; // 35
storage[4388] = -11'b00000100010; // -34
storage[4389] = -11'b00000110101; // -53
storage[4390] = -11'b00000000111; // -7
storage[4391] = -11'b00000011010; // -26
storage[4392] = -11'b00001010111; // -87
storage[4393] = -11'b00000000110; // -6
storage[4394] =  11'b00000000011; // 3
storage[4395] = -11'b00000001000; // -8
storage[4396] = -11'b00010110000; // -176
storage[4397] = -11'b00010111110; // -190
storage[4398] = -11'b00010110101; // -181
storage[4399] =  11'b00000001110; // 14
storage[4400] = -11'b00000000100; // -4
storage[4401] = -11'b00000101010; // -42
storage[4402] =  11'b00000000001; // 1
storage[4403] = -11'b00000001001; // -9
storage[4404] = -11'b00000100011; // -35
storage[4405] = -11'b00000010000; // -16
storage[4406] = -11'b00000111010; // -58
storage[4407] = -11'b00000000101; // -5
storage[4408] =  11'b00000110101; // 53
storage[4409] =  11'b00000111000; // 56
storage[4410] = -11'b00000001100; // -12
storage[4411] =  11'b00000101010; // 42
storage[4412] =  11'b00000011111; // 31
storage[4413] =  11'b00000001011; // 11
storage[4414] = -11'b00000111010; // -58
storage[4415] =  11'b00000000011; // 3
storage[4416] =  11'b00000001110; // 14
storage[4417] = -11'b00000001111; // -15
storage[4418] = -11'b00000000100; // -4
storage[4419] =  11'b00000110010; // 50
storage[4420] = -11'b00000100100; // -36
storage[4421] = -11'b00000100110; // -38
storage[4422] = -11'b00000001110; // -14
storage[4423] =  11'b00000011011; // 27
storage[4424] =  11'b00000110000; // 48
storage[4425] =  11'b00000001111; // 15
storage[4426] =  11'b00001101000; // 104
storage[4427] =  11'b00000100010; // 34
storage[4428] = -11'b00000011111; // -31
storage[4429] =  11'b00000000111; // 7
storage[4430] = -11'b00010000110; // -134
storage[4431] = -11'b00000001100; // -12
storage[4432] = -11'b00000011110; // -30
storage[4433] = -11'b00010111100; // -188
storage[4434] = -11'b00001010011; // -83
storage[4435] =  11'b00001100001; // 97
storage[4436] =  11'b00001010001; // 81
storage[4437] =  11'b00000110100; // 52
storage[4438] =  11'b00000000001; // 1
storage[4439] = -11'b00000100111; // -39
storage[4440] = -11'b00001011010; // -90
storage[4441] = -11'b00000011110; // -30
storage[4442] = -11'b00000011111; // -31
storage[4443] = -11'b00001000110; // -70
storage[4444] =  11'b00001100010; // 98
storage[4445] =  11'b00001010110; // 86
storage[4446] = -11'b00000101011; // -43
storage[4447] = -11'b00000010101; // -21
storage[4448] = -11'b00001011010; // -90
storage[4449] = -11'b00000010111; // -23
storage[4450] =  11'b00000110110; // 54
storage[4451] =  11'b00000001100; // 12
storage[4452] = -11'b00000100101; // -37
storage[4453] =  11'b00000101010; // 42
storage[4454] =  11'b00000110010; // 50
storage[4455] =  11'b00001001001; // 73
storage[4456] =  11'b00000001110; // 14
storage[4457] = -11'b00001001000; // -72
storage[4458] =  11'b00000010010; // 18
storage[4459] = -11'b00000011101; // -29
storage[4460] = -11'b00010101111; // -175
storage[4461] =  11'b00000010101; // 21
storage[4462] = -11'b00010110110; // -182
storage[4463] =  11'b00000101001; // 41
storage[4464] = -11'b00000001010; // -10
storage[4465] =  11'b00000110010; // 50
storage[4466] =  11'b00000101111; // 47
storage[4467] =  11'b00000100110; // 38
storage[4468] =  11'b00000011110; // 30
storage[4469] =  11'b00000000101; // 5
storage[4470] =  11'b00000100000; // 32
storage[4471] =  11'b00000010110; // 22
storage[4472] = -11'b00000101100; // -44
storage[4473] = -11'b00000111111; // -63
storage[4474] = -11'b00000000010; // -2
storage[4475] =  11'b00001010001; // 81
storage[4476] =  11'b00000010010; // 18
storage[4477] = -11'b00000000001; // -1
storage[4478] =  11'b00001001110; // 78
storage[4479] =  11'b00000100011; // 35
storage[4480] =  11'b00001000010; // 66
storage[4481] =  11'b00000010110; // 22
storage[4482] =  11'b00000100101; // 37
storage[4483] =  11'b00000111110; // 62
storage[4484] =  11'b00000011010; // 26
storage[4485] =  11'b00000010000; // 16
storage[4486] =  11'b00000001110; // 14
storage[4487] =  11'b00000001000; // 8
storage[4488] =  11'b00001000110; // 70
storage[4489] = -11'b00000001010; // -10
storage[4490] =  11'b00000100010; // 34
storage[4491] =  11'b00000101000; // 40
storage[4492] =  11'b00000110110; // 54
storage[4493] = -11'b00000000011; // -3
storage[4494] = -11'b00000011000; // -24
storage[4495] =  11'b00000011000; // 24
storage[4496] =  11'b00000001111; // 15
storage[4497] =  11'b00000010000; // 16
storage[4498] = -11'b00000001000; // -8
storage[4499] =  11'b00000000101; // 5
storage[4500] = -11'b00000010010; // -18
storage[4501] =  11'b00001000100; // 68
storage[4502] = -11'b00010000000; // -128
storage[4503] = -11'b00000010000; // -16
storage[4504] =  11'b00001000110; // 70
storage[4505] = -11'b00001100111; // -103
storage[4506] = -11'b00001010001; // -81
storage[4507] =  11'b00000101000; // 40
storage[4508] = -11'b00001111001; // -121
storage[4509] = -11'b00000011011; // -27
storage[4510] = -11'b00000011000; // -24
storage[4511] =  11'b00001001110; // 78
storage[4512] =  11'b00000011011; // 27
storage[4513] = -11'b00000010111; // -23
storage[4514] =  11'b00000110011; // 51
storage[4515] = -11'b00000010011; // -19
storage[4516] = -11'b00011000011; // -195
storage[4517] = -11'b00000110000; // -48
storage[4518] =  11'b00001000101; // 69
storage[4519] =  11'b00000001110; // 14
storage[4520] =  11'b00000100010; // 34
storage[4521] = -11'b00000010001; // -17
storage[4522] = -11'b00000010001; // -17
storage[4523] = -11'b00000000011; // -3
storage[4524] = -11'b00000101111; // -47
storage[4525] =  11'b00001100101; // 101
storage[4526] =  11'b00001000011; // 67
storage[4527] =  11'b00000001010; // 10
storage[4528] = -11'b00000000100; // -4
storage[4529] =  11'b00000110101; // 53
storage[4530] =  11'b00000011110; // 30
storage[4531] = -11'b00001010010; // -82
storage[4532] = -11'b00001101111; // -111
storage[4533] = -11'b00000110100; // -52
storage[4534] =  11'b00000110111; // 55
storage[4535] = -11'b00000100110; // -38
storage[4536] =  11'b00000000100; // 4
storage[4537] = -11'b00000000110; // -6
storage[4538] = -11'b00001011000; // -88
storage[4539] = -11'b00000100110; // -38
storage[4540] = -11'b00000000101; // -5
storage[4541] = -11'b00000010111; // -23
storage[4542] = -11'b00000111110; // -62
storage[4543] =  11'b00000000011; // 3
storage[4544] = -11'b00001010100; // -84
storage[4545] = -11'b00000011100; // -28
storage[4546] =  11'b00000110101; // 53
storage[4547] =  11'b00001001111; // 79
storage[4548] =  11'b00000011100; // 28
storage[4549] =  11'b00000111110; // 62
storage[4550] =  11'b00000000011; // 3
storage[4551] =  11'b00001000101; // 69
storage[4552] = -11'b00000001100; // -12
storage[4553] = -11'b00001000010; // -66
storage[4554] = -11'b00000001111; // -15
storage[4555] =  11'b00000110000; // 48
storage[4556] = -11'b00000000001; // -1
storage[4557] = -11'b00000011100; // -28
storage[4558] =  11'b00000010110; // 22
storage[4559] = -11'b00000000101; // -5
storage[4560] = -11'b00001010001; // -81
storage[4561] =  11'b00000111101; // 61
storage[4562] =  11'b00000111100; // 60
storage[4563] = -11'b00000101101; // -45
storage[4564] = -11'b00001001101; // -77
storage[4565] = -11'b00000100101; // -37
storage[4566] =  11'b00000001001; // 9
storage[4567] =  11'b00000000101; // 5
storage[4568] =  11'b00000000110; // 6
storage[4569] =  11'b00000110111; // 55
storage[4570] =  11'b00000010011; // 19
storage[4571] =  11'b00000110011; // 51
storage[4572] = -11'b00000010101; // -21
storage[4573] =  11'b00000100001; // 33
storage[4574] = -11'b00000000110; // -6
storage[4575] = -11'b00000010110; // -22
storage[4576] = -11'b00001111011; // -123
storage[4577] = -11'b00000100101; // -37
storage[4578] =  11'b00000100100; // 36
storage[4579] = -11'b00010000100; // -132
storage[4580] = -11'b00001011101; // -93
storage[4581] =  11'b00000010101; // 21
storage[4582] =  11'b00000110110; // 54
storage[4583] =  11'b00001001000; // 72
storage[4584] = -11'b00000011100; // -28
storage[4585] =  11'b00000110010; // 50
storage[4586] =  11'b00000100010; // 34
storage[4587] =  11'b00000001001; // 9
storage[4588] =  11'b00000011010; // 26
storage[4589] =  11'b00001001011; // 75
storage[4590] = -11'b00000011110; // -30
storage[4591] =  11'b00000101100; // 44
storage[4592] =  11'b00001000011; // 67
storage[4593] = -11'b00001010011; // -83
storage[4594] =  11'b00001000110; // 70
storage[4595] =  11'b00001010011; // 83
storage[4596] = -11'b00000010101; // -21
storage[4597] =  11'b00001000100; // 68
storage[4598] =  11'b00000001101; // 13
storage[4599] =  11'b00000001100; // 12
storage[4600] = -11'b00000101000; // -40
storage[4601] = -11'b00001001001; // -73
storage[4602] = -11'b00010001011; // -139
storage[4603] = -11'b00000101100; // -44
storage[4604] = -11'b00001110011; // -115
storage[4605] = -11'b00000110100; // -52
storage[4606] = -11'b00001001000; // -72
storage[4607] = -11'b00000010011; // -19
storage[4608] = -11'b00000101000; // -40
storage[4609] = -11'b00000010101; // -21
storage[4610] = -11'b00000101001; // -41
storage[4611] = -11'b00000001110; // -14
storage[4612] =  11'b00000111010; // 58
storage[4613] = -11'b00000001010; // -10
storage[4614] = -11'b00000001100; // -12
storage[4615] =  11'b00000011110; // 30
storage[4616] = -11'b00000011010; // -26
storage[4617] = -11'b00000100000; // -32
storage[4618] = -11'b00000011011; // -27
storage[4619] = -11'b00001000011; // -67
storage[4620] =  11'b00000000101; // 5
storage[4621] =  11'b00000100100; // 36
storage[4622] = -11'b00000000001; // -1
storage[4623] = -11'b00000010011; // -19
storage[4624] =  11'b00000011111; // 31
storage[4625] =  11'b00000111001; // 57
storage[4626] = -11'b00000001001; // -9
storage[4627] = -11'b00000110010; // -50
storage[4628] =  11'b00000010101; // 21
storage[4629] =  11'b00000000111; // 7
storage[4630] = -11'b00010000110; // -134
storage[4631] = -11'b00000111001; // -57
storage[4632] =  11'b00000000010; // 2
storage[4633] = -11'b00000011100; // -28
storage[4634] = -11'b00001100000; // -96
storage[4635] =  11'b00000000100; // 4
storage[4636] = -11'b00000101101; // -45
storage[4637] =  11'b00000101001; // 41
storage[4638] =  11'b00001010000; // 80
storage[4639] = -11'b00000111000; // -56
storage[4640] =  11'b00000111111; // 63
storage[4641] =  11'b00001110110; // 118
storage[4642] = -11'b00000110001; // -49
storage[4643] = -11'b00000000111; // -7
storage[4644] =  11'b00000110011; // 51
storage[4645] = -11'b00000101001; // -41
storage[4646] = -11'b00000100101; // -37
storage[4647] = -11'b00000011001; // -25
storage[4648] = -11'b00000111101; // -61
storage[4649] = -11'b00000010110; // -22
storage[4650] = -11'b00001001100; // -76
storage[4651] =  11'b00000001100; // 12
storage[4652] =  11'b00000001000; // 8
storage[4653] = -11'b00000111011; // -59
storage[4654] =  11'b00000110001; // 49
storage[4655] =  11'b00000001000; // 8
storage[4656] =  11'b00000011100; // 28
storage[4657] = -11'b00001011001; // -89
storage[4658] = -11'b00000111000; // -56
storage[4659] = -11'b00000010000; // -16
storage[4660] = -11'b00000001100; // -12
storage[4661] =  11'b00000011010; // 26
storage[4662] =  11'b00000001001; // 9
storage[4663] = -11'b00000111100; // -60
storage[4664] = -11'b00001010100; // -84
storage[4665] =  11'b00000001101; // 13
storage[4666] = -11'b00000100001; // -33
storage[4667] = -11'b00000001111; // -15
storage[4668] =  11'b00000001110; // 14
storage[4669] = -11'b00000011001; // -25
storage[4670] = -11'b00000001110; // -14
storage[4671] =  11'b00000011001; // 25
storage[4672] = -11'b00000111000; // -56
storage[4673] =  11'b00000001101; // 13
storage[4674] = -11'b00000010001; // -17
storage[4675] = -11'b00001010111; // -87
storage[4676] =  11'b00000000001; // 1
storage[4677] =  11'b00000001011; // 11
storage[4678] =  11'b00000000001; // 1
storage[4679] =  11'b00001100001; // 97
storage[4680] = -11'b00000001001; // -9
storage[4681] = -11'b00000000011; // -3
storage[4682] = -11'b00010011000; // -152
storage[4683] = -11'b00001000011; // -67
storage[4684] = -11'b00000000011; // -3
storage[4685] = -11'b00000010100; // -20
storage[4686] =  11'b00000000101; // 5
storage[4687] = -11'b00000001110; // -14
storage[4688] = -11'b00000100101; // -37
storage[4689] =  11'b00000010000; // 16
storage[4690] = -11'b00001010000; // -80
storage[4691] = -11'b00000010011; // -19
storage[4692] = -11'b00000001111; // -15
storage[4693] = -11'b00001011111; // -95
storage[4694] =  11'b00000010001; // 17
storage[4695] = -11'b00000000010; // -2
storage[4696] = -11'b00000100100; // -36
storage[4697] = -11'b00000010101; // -21
storage[4698] = -11'b00000001001; // -9
storage[4699] =  11'b00000000101; // 5
storage[4700] =  11'b00000001011; // 11
storage[4701] =  11'b00000101110; // 46
storage[4702] =  11'b00000111011; // 59
storage[4703] = -11'b00000011100; // -28
storage[4704] =  11'b00000100101; // 37
storage[4705] =  11'b00001110010; // 114
storage[4706] = -11'b00000100100; // -36
storage[4707] =  11'b00000101100; // 44
storage[4708] =  11'b00000001101; // 13
storage[4709] =  11'b00000101111; // 47
storage[4710] =  11'b00000010111; // 23
storage[4711] =  11'b00000001111; // 15
storage[4712] =  11'b00000011101; // 29
storage[4713] = -11'b00001001010; // -74
storage[4714] =  11'b00000111110; // 62
storage[4715] =  11'b00000101110; // 46
storage[4716] = -11'b00010000111; // -135
storage[4717] = -11'b00000010000; // -16
storage[4718] = -11'b00000000010; // -2
storage[4719] = -11'b00001001111; // -79
storage[4720] = -11'b00000001100; // -12
storage[4721] = -11'b00000010011; // -19
storage[4722] =  11'b00000000000; // 0
storage[4723] = -11'b00001000000; // -64
storage[4724] = -11'b00010111111; // -191
storage[4725] = -11'b00000110001; // -49
storage[4726] = -11'b00000000110; // -6
storage[4727] =  11'b00000011000; // 24
storage[4728] = -11'b00001110101; // -117
storage[4729] = -11'b00000101110; // -46
storage[4730] = -11'b00000100111; // -39
storage[4731] = -11'b00010010011; // -147
storage[4732] = -11'b00001100111; // -103
storage[4733] = -11'b00001100100; // -100
storage[4734] = -11'b00010010011; // -147
storage[4735] =  11'b00001001010; // 74
storage[4736] =  11'b00000110101; // 53
storage[4737] = -11'b00000100011; // -35
storage[4738] = -11'b00000110100; // -52
storage[4739] =  11'b00000110000; // 48
storage[4740] = -11'b00000100100; // -36
storage[4741] = -11'b00000000001; // -1
storage[4742] = -11'b00000011110; // -30
storage[4743] = -11'b00000011100; // -28
storage[4744] =  11'b00001011100; // 92
storage[4745] = -11'b00000101010; // -42
storage[4746] =  11'b00000100001; // 33
storage[4747] =  11'b00000100101; // 37
storage[4748] = -11'b00001000100; // -68
storage[4749] =  11'b00000000001; // 1
storage[4750] =  11'b00000001110; // 14
storage[4751] = -11'b00000001111; // -15
storage[4752] = -11'b00000011001; // -25
storage[4753] = -11'b00000011100; // -28
storage[4754] =  11'b00000001111; // 15
storage[4755] =  11'b00000100000; // 32
storage[4756] =  11'b00000000100; // 4
storage[4757] = -11'b00001000001; // -65
storage[4758] = -11'b00001000101; // -69
storage[4759] =  11'b00001001001; // 73
storage[4760] = -11'b00001010010; // -82
storage[4761] = -11'b00010100000; // -160
storage[4762] =  11'b00001000110; // 70
storage[4763] =  11'b00000111111; // 63
storage[4764] =  11'b00001001001; // 73
storage[4765] =  11'b00000101000; // 40
storage[4766] =  11'b00000101001; // 41
storage[4767] =  11'b00000101110; // 46
storage[4768] =  11'b00000110000; // 48
storage[4769] =  11'b00000100101; // 37
storage[4770] =  11'b00000011001; // 25
storage[4771] = -11'b00000101110; // -46
storage[4772] = -11'b00001000000; // -64
storage[4773] = -11'b00000000001; // -1
storage[4774] =  11'b00000011011; // 27
storage[4775] = -11'b00000101111; // -47
storage[4776] = -11'b00000011101; // -29
storage[4777] =  11'b00000000101; // 5
storage[4778] = -11'b00000010101; // -21
storage[4779] = -11'b00000100100; // -36
storage[4780] =  11'b00001101110; // 110
storage[4781] =  11'b00000111100; // 60
storage[4782] =  11'b00000101111; // 47
storage[4783] = -11'b00001011000; // -88
storage[4784] =  11'b00000001001; // 9
storage[4785] =  11'b00000100110; // 38
storage[4786] = -11'b00000001111; // -15
storage[4787] = -11'b00001010000; // -80
storage[4788] = -11'b00001000011; // -67
storage[4789] = -11'b00000100000; // -32
storage[4790] = -11'b00000100011; // -35
storage[4791] =  11'b00000001111; // 15
storage[4792] = -11'b00010011110; // -158
storage[4793] = -11'b00001110011; // -115
storage[4794] = -11'b00000000110; // -6
storage[4795] = -11'b00001001110; // -78
storage[4796] = -11'b00000010101; // -21
storage[4797] = -11'b00000010101; // -21
storage[4798] = -11'b00000110000; // -48
storage[4799] = -11'b00001111010; // -122
storage[4800] =  11'b00000011101; // 29
storage[4801] =  11'b00000001101; // 13
storage[4802] = -11'b00000110101; // -53
storage[4803] = -11'b00010001001; // -137
storage[4804] =  11'b00000110001; // 49
storage[4805] =  11'b00000010110; // 22
storage[4806] = -11'b00000100100; // -36
storage[4807] = -11'b00000101010; // -42
storage[4808] =  11'b00000101110; // 46
storage[4809] = -11'b00001010001; // -81
storage[4810] = -11'b00000010101; // -21
storage[4811] =  11'b00000000111; // 7
storage[4812] = -11'b00000000100; // -4
storage[4813] =  11'b00000100011; // 35
storage[4814] =  11'b00000011111; // 31
storage[4815] =  11'b00000110101; // 53
storage[4816] = -11'b00000011001; // -25
storage[4817] = -11'b00000001010; // -10
storage[4818] =  11'b00000100000; // 32
storage[4819] =  11'b00000001011; // 11
storage[4820] =  11'b00000010000; // 16
storage[4821] =  11'b00001001011; // 75
storage[4822] =  11'b00000100011; // 35
storage[4823] =  11'b00000000111; // 7
storage[4824] = -11'b00000101100; // -44
storage[4825] =  11'b00000110001; // 49
storage[4826] =  11'b00000101001; // 41
storage[4827] =  11'b00000000100; // 4
storage[4828] =  11'b00000110100; // 52
storage[4829] =  11'b00000010001; // 17
storage[4830] = -11'b00000000100; // -4
storage[4831] = -11'b00000100010; // -34
storage[4832] =  11'b00000110100; // 52
storage[4833] =  11'b00001100011; // 99
storage[4834] =  11'b00000001101; // 13
storage[4835] = -11'b00000010101; // -21
storage[4836] = -11'b00001000011; // -67
storage[4837] = -11'b00000100100; // -36
storage[4838] = -11'b00000010010; // -18
storage[4839] = -11'b00000111111; // -63
storage[4840] =  11'b00000010100; // 20
storage[4841] =  11'b00000000001; // 1
storage[4842] = -11'b00000011110; // -30
storage[4843] =  11'b00000111100; // 60
storage[4844] =  11'b00000111101; // 61
storage[4845] =  11'b00000101101; // 45
storage[4846] = -11'b00000010001; // -17
storage[4847] = -11'b00001000001; // -65
storage[4848] = -11'b00001100000; // -96
storage[4849] =  11'b00000110011; // 51
storage[4850] = -11'b00000101011; // -43
storage[4851] = -11'b00001010001; // -81
storage[4852] =  11'b00000000000; // 0
storage[4853] = -11'b00000100100; // -36
storage[4854] = -11'b00000100010; // -34
storage[4855] =  11'b00000011110; // 30
storage[4856] = -11'b00000001111; // -15
storage[4857] =  11'b00000100011; // 35
storage[4858] = -11'b00000100100; // -36
storage[4859] = -11'b00000010001; // -17
storage[4860] =  11'b00000001101; // 13
storage[4861] =  11'b00000110111; // 55
storage[4862] = -11'b00000111000; // -56
storage[4863] = -11'b00000110000; // -48
storage[4864] = -11'b00001100000; // -96
storage[4865] =  11'b00000000000; // 0
storage[4866] =  11'b00000000100; // 4
storage[4867] = -11'b00001100000; // -96
storage[4868] =  11'b00000111111; // 63
storage[4869] =  11'b00001110010; // 114
storage[4870] =  11'b00000000111; // 7
storage[4871] = -11'b00000010111; // -23
storage[4872] =  11'b00000001001; // 9
storage[4873] = -11'b00000010111; // -23
storage[4874] = -11'b00000101101; // -45
storage[4875] = -11'b00000010111; // -23
storage[4876] =  11'b00000101111; // 47
storage[4877] = -11'b00000100011; // -35
storage[4878] =  11'b00000011000; // 24
storage[4879] = -11'b00000111001; // -57
storage[4880] = -11'b00000010101; // -21
storage[4881] = -11'b00000101100; // -44
storage[4882] = -11'b00000110000; // -48
storage[4883] = -11'b00001010111; // -87
storage[4884] = -11'b00001101000; // -104
storage[4885] = -11'b00000100101; // -37
storage[4886] = -11'b00001110010; // -114
storage[4887] =  11'b00000100000; // 32
storage[4888] =  11'b00001000101; // 69
storage[4889] =  11'b00000111011; // 59
storage[4890] =  11'b00000010101; // 21
storage[4891] =  11'b00001100110; // 102
storage[4892] =  11'b00001011101; // 93
storage[4893] =  11'b00001101110; // 110
storage[4894] = -11'b00000000100; // -4
storage[4895] =  11'b00001010100; // 84
storage[4896] =  11'b00000100001; // 33
storage[4897] =  11'b00000001100; // 12
storage[4898] = -11'b00001000001; // -65
storage[4899] = -11'b00001000010; // -66
storage[4900] = -11'b00001001001; // -73
storage[4901] = -11'b00001001011; // -75
storage[4902] = -11'b00000010101; // -21
storage[4903] = -11'b00000000010; // -2
storage[4904] = -11'b00000101110; // -46
storage[4905] =  11'b00001010011; // 83
storage[4906] = -11'b00000111110; // -62
storage[4907] = -11'b00000001101; // -13
storage[4908] = -11'b00000010000; // -16
storage[4909] =  11'b00000000101; // 5
storage[4910] =  11'b00000101001; // 41
storage[4911] =  11'b00000100011; // 35
storage[4912] = -11'b00000010110; // -22
storage[4913] =  11'b00000001010; // 10
storage[4914] =  11'b00000110110; // 54
storage[4915] = -11'b00000001100; // -12
storage[4916] =  11'b00000001111; // 15
storage[4917] = -11'b00000001010; // -10
storage[4918] =  11'b00000111010; // 58
storage[4919] =  11'b00000011000; // 24
storage[4920] = -11'b00000011111; // -31
storage[4921] = -11'b00001000111; // -71
storage[4922] =  11'b00000010110; // 22
storage[4923] =  11'b00000010011; // 19
storage[4924] =  11'b00001001101; // 77
storage[4925] =  11'b00000011010; // 26
storage[4926] =  11'b00000101000; // 40
storage[4927] = -11'b00000110000; // -48
storage[4928] = -11'b00000000100; // -4
storage[4929] = -11'b00001101100; // -108
storage[4930] = -11'b00000011011; // -27
storage[4931] = -11'b00000010010; // -18
storage[4932] = -11'b00000010111; // -23
storage[4933] = -11'b00000001011; // -11
storage[4934] = -11'b00000010100; // -20
storage[4935] = -11'b00000100111; // -39
storage[4936] =  11'b00001111001; // 121
storage[4937] = -11'b00000001001; // -9
storage[4938] =  11'b00000101110; // 46
storage[4939] = -11'b00000110101; // -53
storage[4940] =  11'b00000001011; // 11
storage[4941] = -11'b00000010011; // -19
storage[4942] =  11'b00000100101; // 37
storage[4943] =  11'b00001001011; // 75
storage[4944] = -11'b00000010001; // -17
storage[4945] = -11'b00000101001; // -41
storage[4946] =  11'b00000001001; // 9
storage[4947] =  11'b00000100100; // 36
storage[4948] = -11'b00001111111; // -127
storage[4949] = -11'b00000001010; // -10
storage[4950] =  11'b00000101000; // 40
storage[4951] = -11'b00000011000; // -24
storage[4952] =  11'b00000011101; // 29
storage[4953] = -11'b00000101011; // -43
storage[4954] =  11'b00000000110; // 6
storage[4955] =  11'b00000100001; // 33
storage[4956] =  11'b00000100010; // 34
storage[4957] = -11'b00001001111; // -79
storage[4958] =  11'b00000111100; // 60
storage[4959] =  11'b00000001101; // 13
storage[4960] = -11'b00001001101; // -77
storage[4961] = -11'b00001000001; // -65
storage[4962] =  11'b00000001000; // 8
storage[4963] = -11'b00001011010; // -90
storage[4964] = -11'b00000100001; // -33
storage[4965] = -11'b00000011101; // -29
storage[4966] = -11'b00000011110; // -30
storage[4967] = -11'b00000011110; // -30
storage[4968] = -11'b00000111001; // -57
storage[4969] = -11'b00000100011; // -35
storage[4970] = -11'b00000001110; // -14
storage[4971] =  11'b00000010111; // 23
storage[4972] =  11'b00000001001; // 9
storage[4973] =  11'b00000110001; // 49
storage[4974] =  11'b00000001111; // 15
storage[4975] =  11'b00001001100; // 76
storage[4976] =  11'b00000111000; // 56
storage[4977] = -11'b00000011101; // -29
storage[4978] =  11'b00000110000; // 48
storage[4979] = -11'b00000001011; // -11
storage[4980] = -11'b00000101000; // -40
storage[4981] =  11'b00000110101; // 53
storage[4982] =  11'b00001001100; // 76
storage[4983] =  11'b00000001000; // 8
storage[4984] = -11'b00000101110; // -46
storage[4985] =  11'b00000001001; // 9
storage[4986] =  11'b00000110000; // 48
storage[4987] =  11'b00001011101; // 93
storage[4988] =  11'b00000110010; // 50
storage[4989] = -11'b00010010010; // -146
storage[4990] =  11'b00000110011; // 51
storage[4991] = -11'b00000000010; // -2
storage[4992] =  11'b00000000010; // 2
storage[4993] =  11'b00000001100; // 12
storage[4994] = -11'b00000010111; // -23
storage[4995] =  11'b00000011100; // 28
storage[4996] =  11'b00000010100; // 20
storage[4997] =  11'b00000001001; // 9
storage[4998] = -11'b00000101111; // -47
storage[4999] =  11'b00000010101; // 21
storage[5000] =  11'b00000101111; // 47
storage[5001] = -11'b00000110000; // -48
storage[5002] =  11'b00000000001; // 1
storage[5003] =  11'b00000001100; // 12
storage[5004] = -11'b00000001111; // -15
storage[5005] =  11'b00000100110; // 38
storage[5006] = -11'b00000000010; // -2
storage[5007] = -11'b00000010100; // -20
storage[5008] = -11'b00000101011; // -43
storage[5009] =  11'b00000100000; // 32
storage[5010] = -11'b00000101111; // -47
storage[5011] = -11'b00000000111; // -7
storage[5012] =  11'b00000000000; // 0
storage[5013] =  11'b00000110100; // 52
storage[5014] =  11'b00000110111; // 55
storage[5015] =  11'b00000110100; // 52
storage[5016] = -11'b00001110100; // -116
storage[5017] =  11'b00000110011; // 51
storage[5018] = -11'b00000011110; // -30
storage[5019] = -11'b00001010011; // -83
storage[5020] =  11'b00001101001; // 105
storage[5021] =  11'b00000011111; // 31
storage[5022] =  11'b00001100010; // 98
storage[5023] =  11'b00001101010; // 106
storage[5024] =  11'b00000011100; // 28
storage[5025] = -11'b00001100110; // -102
storage[5026] = -11'b00000001100; // -12
storage[5027] =  11'b00000111111; // 63
storage[5028] =  11'b00000011000; // 24
storage[5029] =  11'b00000111010; // 58
storage[5030] =  11'b00000000000; // 0
storage[5031] = -11'b00000100001; // -33
storage[5032] = -11'b00000111110; // -62
storage[5033] = -11'b00001011000; // -88
storage[5034] =  11'b00001011001; // 89
storage[5035] =  11'b00000110000; // 48
storage[5036] =  11'b00000011110; // 30
storage[5037] = -11'b00000001110; // -14
storage[5038] =  11'b00000100011; // 35
storage[5039] =  11'b00000010010; // 18
storage[5040] = -11'b00000000010; // -2
storage[5041] =  11'b00000101100; // 44
storage[5042] =  11'b00000010000; // 16
storage[5043] = -11'b00000001001; // -9
storage[5044] = -11'b00000000111; // -7
storage[5045] = -11'b00000010010; // -18
storage[5046] =  11'b00000000110; // 6
storage[5047] =  11'b00000110010; // 50
storage[5048] =  11'b00000110111; // 55
storage[5049] = -11'b00000100000; // -32
storage[5050] =  11'b00010001110; // 142
storage[5051] =  11'b00001000011; // 67
storage[5052] =  11'b00000111000; // 56
storage[5053] =  11'b00000111111; // 63
storage[5054] =  11'b00000000001; // 1
storage[5055] =  11'b00000011011; // 27
storage[5056] =  11'b00000010101; // 21
storage[5057] =  11'b00000001001; // 9
storage[5058] = -11'b00000100001; // -33
storage[5059] = -11'b00000100110; // -38
storage[5060] = -11'b00000100000; // -32
storage[5061] =  11'b00000011001; // 25
storage[5062] = -11'b00001011010; // -90
storage[5063] = -11'b00000100011; // -35
storage[5064] =  11'b00000010001; // 17
storage[5065] = -11'b00001101111; // -111
storage[5066] =  11'b00001000001; // 65
storage[5067] =  11'b00000001000; // 8
storage[5068] =  11'b00000110001; // 49
storage[5069] =  11'b00000100110; // 38
storage[5070] =  11'b00000001011; // 11
storage[5071] = -11'b00001000111; // -71
storage[5072] = -11'b00000001111; // -15
storage[5073] =  11'b00001000010; // 66
storage[5074] = -11'b00000101101; // -45
storage[5075] = -11'b00000111000; // -56
storage[5076] =  11'b00000110111; // 55
storage[5077] =  11'b00000110110; // 54
storage[5078] = -11'b00000010110; // -22
storage[5079] = -11'b00000001000; // -8
storage[5080] = -11'b00001000011; // -67
storage[5081] =  11'b00000010010; // 18
storage[5082] =  11'b00000011110; // 30
storage[5083] =  11'b00000010010; // 18
storage[5084] = -11'b00000000001; // -1
storage[5085] = -11'b00000010011; // -19
storage[5086] =  11'b00000001011; // 11
storage[5087] = -11'b00000010101; // -21
storage[5088] = -11'b00000101001; // -41
storage[5089] =  11'b00000100101; // 37
storage[5090] = -11'b00000010011; // -19
storage[5091] = -11'b00000010100; // -20
storage[5092] = -11'b00000101001; // -41
storage[5093] =  11'b00000011110; // 30
storage[5094] =  11'b00000110000; // 48
storage[5095] = -11'b00001111111; // -127
storage[5096] = -11'b00000001010; // -10
storage[5097] = -11'b00000001000; // -8
storage[5098] = -11'b00000100100; // -36
storage[5099] =  11'b00001011100; // 92
storage[5100] =  11'b00000001001; // 9
storage[5101] = -11'b00000001011; // -11
storage[5102] =  11'b00000101001; // 41
storage[5103] =  11'b00000011110; // 30
storage[5104] = -11'b00000110100; // -52
storage[5105] = -11'b00000000100; // -4
storage[5106] = -11'b00001000101; // -69
storage[5107] = -11'b00000111110; // -62
storage[5108] = -11'b00000111000; // -56
storage[5109] = -11'b00000110010; // -50
storage[5110] =  11'b00000000000; // 0
storage[5111] =  11'b00000010111; // 23
storage[5112] =  11'b00000100010; // 34
storage[5113] =  11'b00000010010; // 18
storage[5114] = -11'b00000011000; // -24
storage[5115] = -11'b00000011111; // -31
storage[5116] = -11'b00001000100; // -68
storage[5117] = -11'b00000111111; // -63
storage[5118] = -11'b00000110000; // -48
storage[5119] = -11'b00000011011; // -27
storage[5120] = -11'b00001000111; // -71
storage[5121] = -11'b00001000100; // -68
storage[5122] =  11'b00000110011; // 51
storage[5123] =  11'b00000100100; // 36
storage[5124] =  11'b00000101001; // 41
storage[5125] =  11'b00000100011; // 35
storage[5126] =  11'b00000111111; // 63
storage[5127] =  11'b00000011000; // 24
storage[5128] =  11'b00000000100; // 4
storage[5129] = -11'b00000001111; // -15
storage[5130] = -11'b00000100011; // -35
storage[5131] = -11'b00000010101; // -21
storage[5132] = -11'b00000111100; // -60
storage[5133] = -11'b00010011001; // -153
storage[5134] =  11'b00000000111; // 7
storage[5135] = -11'b00000011101; // -29
storage[5136] = -11'b00010010000; // -144
storage[5137] =  11'b00000111001; // 57
storage[5138] =  11'b00000011100; // 28
storage[5139] = -11'b00000100101; // -37
storage[5140] =  11'b00000010100; // 20
storage[5141] =  11'b00000000100; // 4
storage[5142] =  11'b00001010010; // 82
storage[5143] = -11'b00000000100; // -4
storage[5144] =  11'b00000010111; // 23
storage[5145] =  11'b00001000000; // 64
storage[5146] =  11'b00000011110; // 30
storage[5147] =  11'b00000011001; // 25
storage[5148] = -11'b00000110101; // -53
storage[5149] = -11'b00001100011; // -99
storage[5150] = -11'b00000111011; // -59
storage[5151] = -11'b00000111101; // -61
storage[5152] = -11'b00001011001; // -89
storage[5153] = -11'b00010110101; // -181
storage[5154] = -11'b00000010000; // -16
storage[5155] = -11'b00001000101; // -69
storage[5156] = -11'b00001000111; // -71
storage[5157] =  11'b00000011110; // 30
storage[5158] = -11'b00000100100; // -36
storage[5159] = -11'b00001100001; // -97
storage[5160] = -11'b00000110001; // -49
storage[5161] =  11'b00000001010; // 10
storage[5162] = -11'b00000001010; // -10
storage[5163] =  11'b00000001111; // 15
storage[5164] = -11'b00010001010; // -138
storage[5165] = -11'b00001100111; // -103
storage[5166] = -11'b00001000110; // -70
storage[5167] =  11'b00001010011; // 83
storage[5168] =  11'b00001111000; // 120
storage[5169] =  11'b00000100111; // 39
storage[5170] =  11'b00000011011; // 27
storage[5171] =  11'b00001100000; // 96
storage[5172] =  11'b00000111110; // 62
storage[5173] = -11'b00001000010; // -66
storage[5174] = -11'b00001010111; // -87
storage[5175] = -11'b00001001001; // -73
storage[5176] = -11'b00000100010; // -34
storage[5177] = -11'b00001100010; // -98
storage[5178] = -11'b00000001100; // -12
storage[5179] = -11'b00000000001; // -1
storage[5180] = -11'b00000100111; // -39
storage[5181] =  11'b00000000101; // 5
storage[5182] =  11'b00000111100; // 60
storage[5183] = -11'b00000000001; // -1
storage[5184] = -11'b00000110001; // -49
storage[5185] =  11'b00000010011; // 19
storage[5186] = -11'b00000000111; // -7
storage[5187] =  11'b00000000110; // 6
storage[5188] =  11'b00000010001; // 17
storage[5189] =  11'b00000001000; // 8
storage[5190] = -11'b00000101101; // -45
storage[5191] =  11'b00000011010; // 26
storage[5192] = -11'b00000010010; // -18
storage[5193] = -11'b00000111101; // -61
storage[5194] = -11'b00000011001; // -25
storage[5195] = -11'b00010001111; // -143
storage[5196] =  11'b00000001101; // 13
storage[5197] = -11'b00000000101; // -5
storage[5198] = -11'b00000100001; // -33
storage[5199] = -11'b00000000001; // -1
storage[5200] = -11'b00000111011; // -59
storage[5201] = -11'b00001100110; // -102
storage[5202] = -11'b00000011000; // -24
storage[5203] = -11'b00011110010; // -242
storage[5204] = -11'b00011000000; // -192
storage[5205] = -11'b00000001110; // -14
storage[5206] =  11'b00000001011; // 11
storage[5207] = -11'b00011001010; // -202
storage[5208] = -11'b00010011010; // -154
storage[5209] =  11'b00000101011; // 43
storage[5210] = -11'b00010001001; // -137
storage[5211] = -11'b00010100000; // -160
storage[5212] =  11'b00001010000; // 80
storage[5213] = -11'b00000101001; // -41
storage[5214] =  11'b00000000000; // 0
storage[5215] = -11'b00000110110; // -54
storage[5216] = -11'b00000110100; // -52
storage[5217] =  11'b00000010110; // 22
storage[5218] = -11'b00001101001; // -105
storage[5219] = -11'b00001001011; // -75
storage[5220] =  11'b00000101010; // 42
storage[5221] = -11'b00000110000; // -48
storage[5222] =  11'b00000010010; // 18
storage[5223] = -11'b00010101101; // -173
storage[5224] = -11'b00000001100; // -12
storage[5225] = -11'b00001100001; // -97
storage[5226] = -11'b00000010010; // -18
storage[5227] = -11'b00001010110; // -86
storage[5228] = -11'b00001011110; // -94
storage[5229] = -11'b00000101101; // -45
storage[5230] = -11'b00000000101; // -5
storage[5231] =  11'b00000101010; // 42
storage[5232] = -11'b00000000101; // -5
storage[5233] = -11'b00000000100; // -4
storage[5234] = -11'b00000101011; // -43
storage[5235] = -11'b00000110101; // -53
storage[5236] =  11'b00000111000; // 56
storage[5237] = -11'b00000100101; // -37
storage[5238] = -11'b00000111010; // -58
storage[5239] =  11'b00001100101; // 101
storage[5240] =  11'b00000100101; // 37
storage[5241] = -11'b00000000111; // -7
storage[5242] =  11'b00001001110; // 78
storage[5243] =  11'b00000001101; // 13
storage[5244] =  11'b00001000010; // 66
storage[5245] =  11'b00000011010; // 26
storage[5246] =  11'b00000001101; // 13
storage[5247] = -11'b00000010011; // -19
storage[5248] =  11'b00001010110; // 86
storage[5249] =  11'b00000111010; // 58
storage[5250] = -11'b00000011100; // -28
storage[5251] =  11'b00000111111; // 63
storage[5252] =  11'b00000100000; // 32
storage[5253] = -11'b00000111110; // -62
storage[5254] = -11'b00000100111; // -39
storage[5255] = -11'b00000011101; // -29
storage[5256] = -11'b00011000011; // -195
storage[5257] = -11'b00000000111; // -7
storage[5258] =  11'b00000101010; // 42
storage[5259] = -11'b00000110100; // -52
storage[5260] =  11'b00000011111; // 31
storage[5261] = -11'b00000000010; // -2
storage[5262] =  11'b00000010100; // 20
storage[5263] =  11'b00000111001; // 57
storage[5264] =  11'b00000101011; // 43
storage[5265] =  11'b00000110001; // 49
storage[5266] = -11'b00000101100; // -44
storage[5267] = -11'b00000000001; // -1
storage[5268] =  11'b00000011011; // 27
storage[5269] =  11'b00000010110; // 22
storage[5270] =  11'b00000111010; // 58
storage[5271] =  11'b00000001101; // 13
storage[5272] =  11'b00001100000; // 96
storage[5273] =  11'b00001000000; // 64
storage[5274] =  11'b00001000101; // 69
storage[5275] = -11'b00000001101; // -13
storage[5276] =  11'b00000101100; // 44
storage[5277] =  11'b00001100111; // 103
storage[5278] =  11'b00000000101; // 5
storage[5279] =  11'b00000101100; // 44
storage[5280] =  11'b00000011110; // 30
storage[5281] =  11'b00000011001; // 25
storage[5282] = -11'b00000001010; // -10
storage[5283] = -11'b00000010111; // -23
storage[5284] = -11'b00010010000; // -144
storage[5285] = -11'b00011100101; // -229
storage[5286] = -11'b00001110001; // -113
storage[5287] = -11'b00001001111; // -79
storage[5288] = -11'b00001101001; // -105
storage[5289] = -11'b00001110100; // -116
storage[5290] = -11'b00000010000; // -16
storage[5291] =  11'b00010101101; // 173
storage[5292] = -11'b00010011001; // -153
storage[5293] =  11'b00011000100; // 196
storage[5294] =  11'b00011010011; // 211
storage[5295] =  11'b00000100010; // 34
storage[5296] = -11'b00001010101; // -85
storage[5297] =  11'b00001010100; // 84
storage[5298] = -11'b00010001101; // -141
storage[5299] =  11'b00011000000; // 192
storage[5300] = -11'b00001010001; // -81
storage[5301] = -11'b00000000111; // -7
storage[5302] =  11'b00010100110; // 166
storage[5303] = -11'b00010111001; // -185
storage[5304] =  11'b00000111000; // 56
storage[5305] = -11'b00001001100; // -76
storage[5306] = -11'b00000011110; // -30
storage[5307] = -11'b00000110011; // -51
storage[5308] =  11'b00011101000; // 232
storage[5309] = -11'b00000011010; // -26
storage[5310] = -11'b00010110101; // -181
storage[5311] =  11'b00001101000; // 104
storage[5312] = -11'b00011001111; // -207
storage[5313] =  11'b00001000010; // 66
storage[5314] =  11'b00100000010; // 258
storage[5315] = -11'b00000011011; // -27
storage[5316] = -11'b00011011010; // -218
storage[5317] =  11'b00100100010; // 290
storage[5318] =  11'b00010001001; // 137
storage[5319] = -11'b00010100001; // -161
storage[5320] =  11'b00001000000; // 64
storage[5321] =  11'b00000000001; // 1
storage[5322] =  11'b00001000011; // 67
storage[5323] = -11'b00000100110; // -38
storage[5324] = -11'b00000100000; // -32
storage[5325] = -11'b00000001110; // -14
storage[5326] =  11'b00000100011; // 35
storage[5327] =  11'b00010001011; // 139
storage[5328] = -11'b00101000011; // -323
storage[5329] = -11'b00000100011; // -35
storage[5330] = -11'b00000001100; // -12
storage[5331] = -11'b00010000000; // -128
storage[5332] =  11'b00001010100; // 84
storage[5333] = -11'b00010000100; // -132
storage[5334] =  11'b00011001010; // 202
storage[5335] =  11'b00001001000; // 72
storage[5336] = -11'b00010001110; // -142
storage[5337] =  11'b00000010110; // 22
storage[5338] =  11'b00001111001; // 121
storage[5339] = -11'b00001110111; // -119
storage[5340] = -11'b00010010011; // -147
storage[5341] = -11'b00010011000; // -152
storage[5342] = -11'b00010000000; // -128
storage[5343] =  11'b00000101110; // 46
storage[5344] =  11'b00100001110; // 270
storage[5345] =  11'b00001100011; // 99
storage[5346] =  11'b00000101100; // 44
storage[5347] = -11'b00000101011; // -43
storage[5348] = -11'b00100010110; // -278
storage[5349] =  11'b00001001110; // 78
storage[5350] =  11'b00000111001; // 57
storage[5351] =  11'b00001111110; // 126
storage[5352] = -11'b00010111001; // -185
storage[5353] = -11'b00010000001; // -129
storage[5354] = -11'b00001011111; // -95
storage[5355] = -11'b00000100111; // -39
storage[5356] = -11'b00000110010; // -50
storage[5357] =  11'b00100001011; // 267
storage[5358] = -11'b00010110000; // -176
storage[5359] =  11'b00001000110; // 70
storage[5360] = -11'b00001010011; // -83
storage[5361] =  11'b00010111101; // 189
storage[5362] = -11'b00000011011; // -27
storage[5363] = -11'b00000001100; // -12
storage[5364] =  11'b00000001000; // 8
storage[5365] = -11'b00000100100; // -36
storage[5366] = -11'b00001010101; // -85
storage[5367] = -11'b00011001110; // -206
storage[5368] =  11'b00001000000; // 64
storage[5369] = -11'b00010101011; // -171
storage[5370] = -11'b00000010011; // -19
storage[5371] = -11'b00000011000; // -24
storage[5372] = -11'b00011011101; // -221
storage[5373] =  11'b00000101011; // 43
storage[5374] =  11'b00010011001; // 153
storage[5375] =  11'b00001011110; // 94
storage[5376] = -11'b00011000010; // -194
storage[5377] =  11'b00001101101; // 109
storage[5378] =  11'b00100100011; // 291
storage[5379] = -11'b00010010110; // -150
storage[5380] =  11'b00100000101; // 261
storage[5381] =  11'b00011101011; // 235
storage[5382] = -11'b00100101101; // -301
storage[5383] = -11'b00000010001; // -17
storage[5384] = -11'b00100010101; // -277
storage[5385] = -11'b00000110110; // -54
storage[5386] = -11'b00101011001; // -345
storage[5387] = -11'b00001010000; // -80
storage[5388] = -11'b00011000000; // -192
storage[5389] =  11'b00001001010; // 74
storage[5390] = -11'b00000101100; // -44
storage[5391] = -11'b00011010101; // -213
storage[5392] =  11'b00001100010; // 98
storage[5393] = -11'b00011111001; // -249
storage[5394] = -11'b00001101101; // -109
storage[5395] =  11'b00100110000; // 304
storage[5396] = -11'b00011011100; // -220
storage[5397] =  11'b00010011001; // 153
storage[5398] =  11'b00011110101; // 245
storage[5399] = -11'b00001000000; // -64
storage[5400] = -11'b00001101011; // -107
storage[5401] =  11'b00010000010; // 130
storage[5402] =  11'b00100100111; // 295
storage[5403] = -11'b00011111001; // -249
storage[5404] =  11'b00001110110; // 118
storage[5405] =  11'b00000011011; // 27
storage[5406] =  11'b00001010111; // 87
storage[5407] = -11'b00101010001; // -337
storage[5408] = -11'b00011101101; // -237
storage[5409] = -11'b00000111100; // -60
storage[5410] = -11'b00000100011; // -35
storage[5411] = -11'b00010110000; // -176
storage[5412] = -11'b00010001101; // -141
storage[5413] =  11'b00010010001; // 145
storage[5414] = -11'b00100100110; // -294
storage[5415] =  11'b00010010111; // 151
storage[5416] =  11'b00011111101; // 253
storage[5417] = -11'b00001100101; // -101
storage[5418] = -11'b00011100101; // -229
storage[5419] =  11'b00100011110; // 286
storage[5420] = -11'b00100100010; // -290
storage[5421] = -11'b00010100110; // -166
storage[5422] = -11'b00000100001; // -33
storage[5423] = -11'b00111010101; // -469
storage[5424] = -11'b00001010010; // -82
storage[5425] =  11'b00010010110; // 150
storage[5426] = -11'b00010001010; // -138
storage[5427] =  11'b00010100110; // 166
storage[5428] =  11'b00010010000; // 144
storage[5429] =  11'b00011010100; // 212
storage[5430] = -11'b00100110011; // -307
storage[5431] = -11'b00011010000; // -208
storage[5432] = -11'b00010010111; // -151
storage[5433] = -11'b00100100101; // -293
storage[5434] = -11'b00001111110; // -126
storage[5435] =  11'b00100000000; // 256
storage[5436] =  11'b00001100111; // 103
storage[5437] = -11'b00010010001; // -145
storage[5438] = -11'b00000101010; // -42
storage[5439] = -11'b00010101001; // -169
storage[5440] =  11'b00010000101; // 133
storage[5441] = -11'b00001011000; // -88
storage[5442] =  11'b00001000011; // 67
storage[5443] =  11'b00001110001; // 113
storage[5444] =  11'b01001001010; // 586
storage[5445] =  11'b00011001001; // 201
storage[5446] = -11'b01000111101; // -573
storage[5447] = -11'b01011000010; // -706
storage[5448] = -11'b01010101001; // -681
storage[5449] =  11'b01000000101; // 517
storage[5450] =  11'b00001010011; // 83
storage[5451] =  11'b00000110101; // 53
storage[5452] = -11'b01010010001; // -657
storage[5453] = -11'b00011101011; // -235
storage[5454] = -11'b01110100011; // -931
storage[5455] =  11'b00001011110; // 94
storage[5456] = -11'b00000101011; // -43
storage[5457] =  11'b01010100110; // 678
storage[5458] = -11'b01000011000; // -536
storage[5459] =  11'b00110110001; // 433
end

always @(posedge clk) if (we==1) storage[address_p] <= dp;
always @(posedge clk) if (re==1) datata<=storage[address];

endmodule
